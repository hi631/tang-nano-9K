//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Fri Nov 25 17:18:09 2022

module Gowin_pROM_bios (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hE7E6E6E633B0018EFC646520320A6153006369206F2032284950532D4E54314E;
defparam prom_inst_0.INIT_RAM_01 = 256'h54F7C74C01C74469C72404C71C44A58B028D04076A3C754000F48033F0C0E715;
defparam prom_inst_0.INIT_RAM_02 = 256'hA7AE00000B84003E8384630F1E1E02C7C6440480F6076AD090C7684AC760E0C7;
defparam prom_inst_0.INIT_RAM_03 = 256'hE68710E6746CAA13E315E873646400C6B207E875A8ABE8CE23F8E81913FF1319;
defparam prom_inst_0.INIT_RAM_04 = 256'h65732019DBB8E3E8061076BE00133DE894E813000006021403E7A170B88AB00C;
defparam prom_inst_0.INIT_RAM_05 = 256'h8906B03C07C07524088B50300D3668202020527374334D2C4D20383820430A74;
defparam prom_inst_0.INIT_RAM_06 = 256'h01F580BF078AC540759617E4061FCDCDA8FEA8B4CDC6470700137F57831F1E1F;
defparam prom_inst_0.INIT_RAM_07 = 256'h741E31CA08C90275EB0551803CE2AA027575FFEA720F0CE418E1803CC9E0E9CD;
defparam prom_inst_0.INIT_RAM_08 = 256'h0AF6C0001AA106108AC25B5254E85CE2FBE10275EB81CA80C11DE98486F7EBF7;
defparam prom_inst_0.INIT_RAM_09 = 256'h740404F302F63CF34077B3C2D7BB1A756C148A590EB9BF088AC25B5200802075;
defparam prom_inst_0.INIT_RAM_0A = 256'hC177168056C37580E6E6F81F0E16E8B40CC507048AF716C8EB0A2648F8870398;
defparam prom_inst_0.INIT_RAM_0B = 256'hB774008087EBB4EB868D026BB1E609F401CF00AB76F3E65100372401055EFFE6;
defparam prom_inst_0.INIT_RAM_0C = 256'h50D0D060F0B00007FF00616D656308590246539D072C586CFF078A8350B3EB81;
defparam prom_inst_0.INIT_RAM_0D = 256'h0001BF6975EB6900C74AB4190097C70700BB4C50C74200B60640B8EF00B2B8B8;
defparam prom_inst_0.INIT_RAM_0E = 256'hE880000000060001BF031E008F00C74AB43CEFEF03A0060001BF3C28F9064006;
defparam prom_inst_0.INIT_RAM_0F = 256'h10B9CD10B8EE6FC4B058BA3C96FFF3967506CDABB9C018EFEF8AB0D450403C50;
defparam prom_inst_0.INIT_RAM_10 = 256'hC15BB0B00303C65262753E89078A588A8AD4C910F6896100B0C0B00E8BDBB800;
defparam prom_inst_0.INIT_RAM_11 = 256'h00FF0700CA06EFEF8A00E0E3C18B02400213B8B4B48AB83C3C008AFC000050E3;
defparam prom_inst_0.INIT_RAM_12 = 256'hFF8A5003C0C050EB87E35B0400C35050868AF706036007FEF3B0F3FAA58A7274;
defparam prom_inst_0.INIT_RAM_13 = 256'hB7FE84FEEBEB01EB733A0074747474F800C31000B45003625359C3FF5358FBFB;
defparam prom_inst_0.INIT_RAM_14 = 256'h0061EEC0DACA2E8B3C7B696969FFE9696969E669697A6A3E260600EBCD000006;
defparam prom_inst_0.INIT_RAM_15 = 256'h5AEEC4038AC361F3808AB08B584AC3BABA613089E0A23232E6EEC0DA61FE0F0F;
defparam prom_inst_0.INIT_RAM_16 = 256'h1493BA5AC6C30342C7608AECE042BA50C7B0030C106FD0026F84EC60266B038B;
defparam prom_inst_0.INIT_RAM_17 = 256'h0311C7C7A03EA2011F74F6595103E992D9C310EED66B978A08CD8AC303C0E62E;
defparam prom_inst_0.INIT_RAM_18 = 256'h017400000101DE1EC37C8E611006002E00EB8BBB747674743CA8A8A8A86F5803;
defparam prom_inst_0.INIT_RAM_19 = 256'h89F6FB03838AFBC8DCBA0E8B088BFF0C72C40E808A8B10BD21BD3C07B9614800;
defparam prom_inst_0.INIT_RAM_1A = 256'h743EB874140200F312498CB84700747761B4A8E88B898A742609FFEE6000B030;
defparam prom_inst_0.INIT_RAM_1B = 256'hA11E4F2525250A0C12252574278E7B2600EF000DC4F3B1ABE8A024AB93BB0003;
defparam prom_inst_0.INIT_RAM_1C = 256'hEFEFEFEFEEEFEFEFEEEECFF6088B00001FFFFEED14140880108074366A1F1FCF;
defparam prom_inst_0.INIT_RAM_1D = 256'hF7D500007404807437F6EBC38AE98001DF0880E2C1748B8BFAEFEFEFEEEEEFEE;
defparam prom_inst_0.INIT_RAM_1E = 256'hB48003BD3233C80686033D3EDA830A8B000780988000C3C13ECA8308ECC58C03;
defparam prom_inst_0.INIT_RAM_1F = 256'h1F52B458448912E8648900C700C703C74404088B50FA041A442BFF548B025F8B;
defparam prom_inst_0.INIT_RAM_20 = 256'hFF75FB7452EEC2208AE08A5A321F428AC2037405804A8A1F744E0DC142ECC2F6;
defparam prom_inst_0.INIT_RAM_21 = 256'h91C8838B3BDBDB0000E8B5E81A7C8A1C1F00A21716600000F402C00CFF0C33F8;
defparam prom_inst_0.INIT_RAM_22 = 256'h8665C2090C116B881D29838034803807A2F02EEFBCE8FF850B7473D174F7A4C8;
defparam prom_inst_0.INIT_RAM_23 = 256'h1F87EF9C0375066AEB07A8B85B0707DB6A531FCD889E9C839A98E72226014000;
defparam prom_inst_0.INIT_RAM_24 = 256'h02CBFAB4A7EB028068AA03F6E46772E0E702EB8C893C72743C7258B010503C8A;
defparam prom_inst_0.INIT_RAM_25 = 256'h3C3C727440A81F1E44FC6414E79A805A988BE87297E81FA5A2F672B3E8E953FF;
defparam prom_inst_0.INIT_RAM_26 = 256'h8052FC000A00840400EB36000136004600005E1C1AEB898B8200FACDCFB03C3C;
defparam prom_inst_0.INIT_RAM_27 = 256'h7588DCE80100D842F0E6B8E8077324FB3897B7C000013272185BDBB40E00B4DF;
defparam prom_inst_0.INIT_RAM_28 = 256'h70700E1612801E00057C00BA020A2E30302C30313252207420626165656F6F01;
defparam prom_inst_0.INIT_RAM_29 = 256'h5CACACFB44A33E21069C0300678BB41E1FC0809800C600032E01F61E0000001F;
defparam prom_inst_0.INIT_RAM_2A = 256'h3CDCFF1A2073240A64035A8AB08473240B6403C3E4E481D0EC424202FADACF08;
defparam prom_inst_0.INIT_RAM_2B = 256'hE8DFC3E9EDD1909001C3CD0AB45A30F1C036330026B1F68384BB8906C3B000C3;
defparam prom_inst_0.INIT_RAM_2C = 256'h29800F8E8CC74106C044E9FBB4F40183C2F5F6F580FF3300BBDB472ADBC00265;
defparam prom_inst_0.INIT_RAM_2D = 256'hEAFEB0FD0F8E8CC6CADD064C44E9B4F40183C2C3FFC0EB05FF0E1183034FE8FF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFEF763E8EBAA581FE166FED3CCE8CDB49BB9571EF9FEB3E874C673C704E4E8FE;
defparam prom_inst_0.INIT_RAM_2F = 256'h2A0000FF0000FF0000870000C38BFEC041F63FFC12FE7EE4E8D958FE162B95BE;
defparam prom_inst_0.INIT_RAM_30 = 256'h3F3F00003F2F002F3F003F322D28201C18110E0B05003F3F15153F152A2A0000;
defparam prom_inst_0.INIT_RAM_31 = 256'h3F152A2A00002A002A2A00002A000D0905013F371F373F1F003F3F00103F1000;
defparam prom_inst_0.INIT_RAM_32 = 256'h15153F153F3F15153F152A2A00002A002A2A00002A003F3F15153F153F3F1515;
defparam prom_inst_0.INIT_RAM_33 = 256'h2A002A3F15003F152A2A15002A152A3F00003F002A2A00002A00151105013F3F;
defparam prom_inst_0.INIT_RAM_34 = 256'h1205443933523D3905013F3F15153F153F2A15152A153F3F00153F003F2A0015;
defparam prom_inst_0.INIT_RAM_35 = 256'h016113731A7A11710000504B3F4D473500232124005A27353E0E0730160B001A;
defparam prom_inst_0.INIT_RAM_36 = 256'h0A6A0D6D19790767086802620E6E127214740666167605650464187803631777;
defparam prom_inst_0.INIT_RAM_37 = 256'h000000000000000000000000000000000000000010700C6C0F6F09690B6B1575;
defparam prom_inst_0.INIT_RAM_38 = 256'h0033003400320031006000090000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h003D1B5B00271F2D003B002F002F002E00390030002C003800371E3600352020;
defparam prom_inst_0.INIT_RAM_3A = 256'h002B00001B1B0000000000000000000000000000000000007F081C5C1D5D0A0D;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000002A002D0000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h3930F0EA00000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h06216140C0366AD0B80D6364200072444D6874446C4E30434F436F3961613865;
defparam prom_inst_1.INIT_RAM_01 = 256'h00EF0600EE0600E50600E30600083344B9F50033001602423314F3FF1F078CB8;
defparam prom_inst_1.INIT_RAM_02 = 256'hE6E6CD10C68940C78480D40EC78383444408F8F333334001F40600F40600F206;
defparam prom_inst_1.INIT_RAM_03 = 256'h641300640913757210B199FBE8B0B00613B4B90E1375AF13B43CBF4972F8E200;
defparam prom_inst_1.INIT_RAM_04 = 256'h74654D50CD050069BE00134A10F6E0700091BEE00E1572D03301E6E600C46003;
defparam prom_inst_1.INIT_RAM_05 = 256'h46408006251AF7F88AEC533A0A627A37443141292032682049284D3638500065;
defparam prom_inst_1.INIT_RAM_06 = 256'hB410F511B3E510741F0000606ACF097420CC01041C4702007581020207BB535B;
defparam prom_inst_1.INIT_RAM_07 = 256'h08F63C08EB08741348803CCA36FD75EB0524F6000001740C8A3CC9E10275C815;
defparam prom_inst_1.INIT_RAM_08 = 256'hF6C1E9CD00807175D30472E8BB08BBFBEBFB741373CA04C9027507C006FD0480;
defparam prom_inst_1.INIT_RAM_09 = 256'h02F67402B3C22502740A02033367E4E2F6A84575070CC0E9D30472E8BB527505;
defparam prom_inst_1.INIT_RAM_0A = 256'hEE0E80FC6AFB02FF320A75619617EAED40587432C28059B40BA219780AD8D8C1;
defparam prom_inst_1.INIT_RAM_0B = 256'h0006808A00C900D1E08702C377F30051B481B05F332EB95701743C72741F94FE;
defparam prom_inst_1.INIT_RAM_0C = 256'hBA0E1606800A004099016369206F00E600E641CB920A9D0F750492E052E5ADC3;
defparam prom_inst_1.INIT_RAM_0D = 256'h50C72800193F0020060011BF3CF906BF4000000006B8E6E677EF07B0EFCE0402;
defparam prom_inst_1.INIT_RAM_0E = 256'hA233A0F7C74C50C750E93CF7C7000600412658B8B8504C50C728245D3C69EB4C;
defparam prom_inst_1.INIT_RAM_0F = 256'hF60710B814B0E6EE10BADA0840A0AB33168710B808BFFF58B8E012031E800351;
defparam prom_inst_1.INIT_RAM_10 = 256'hEB580E0F50C26B33001E495783C7C3E1E503FE74060EC3CD1300020716B91208;
defparam prom_inst_1.INIT_RAM_11 = 256'h910302684187618AE3BA028BEBA1B03CC7B8000203400A0313A0F80CC35B8B0E;
defparam prom_inst_1.INIT_RAM_12 = 256'h1EE306DB50868E070000C300C3692A03C6D8DE00CA0661CFAB2002FE03C80F13;
defparam prom_inst_1.INIT_RAM_13 = 256'h07CE00C6F0F480FC1016CD1822181A5108F75AB40AC1DB00525B028851C359F3;
defparam prom_inst_1.INIT_RAM_14 = 256'h8BC38A0303C3FFF01BEBEBEAEAEAEAEAEAEAEAEAEAEAEA624A4924CC104A8A8A;
defparam prom_inst_1.INIT_RAM_15 = 256'h588AEEEEC350C3B0FBC707FA5AEEEEC0DAC30600026FC3C3C02E0303C3CBCD26;
defparam prom_inst_1.INIT_RAM_16 = 256'hE85AC6C30352F342038BF48AEC42C752EE14C002EEE6D8C0E6DBBABA6EC993F2;
defparam prom_inst_1.INIT_RAM_17 = 256'hEC50A80C6F8584F650316140F38B108761FECD8A03C900D56B10F9E3C0EB808A;
defparam prom_inst_1.INIT_RAM_18 = 256'h890313801F8C8933608CDEC3CD0E01DF10092E007A60373020EBEDEEEFE6EEB0;
defparam prom_inst_1.INIT_RAM_19 = 256'h00D83100E10E1000000007AC03F30701182E6AFF160E0700CD0023BD08C3A299;
defparam prom_inst_1.INIT_RAM_1A = 256'h0D49000FBBB0ABA4B900C8AEED2E030CC302018FFC545E058A5074088BC31206;
defparam prom_inst_1.INIT_RAM_1B = 256'h106AEDE8E8E8EDECEAE8E8E9E9E8E8E8000C0400C3AB06B004872FA0AB080D80;
defparam prom_inst_1.INIT_RAM_1C = 256'h252525F425DB3425D1DBC9DCD0EC0880889601078BB4B4FC80FC139240CFA11E;
defparam prom_inst_1.INIT_RAM_1D = 256'hD959595018F675E7F6EB08BD26B47500B4EB360AE91FD10E80A7F46B7525F4C9;
defparam prom_inst_1.INIT_RAM_1E = 256'h06FABDB2F6C0BA0CC4B8FEF700E8C1D0A175FAB4FA008383F749E16B068AD88E;
defparam prom_inst_1.INIT_RAM_1F = 256'h8B5601B4186C89061044894489448944021A33ECA18007E40244D50A44C41ADC;
defparam prom_inst_1.INIT_RAM_20 = 256'h0125ECFBEC5AFB74E0EBE042C0EE8AC4FDD305B8EE4AC8CF33744EEE4224038B;
defparam prom_inst_1.INIT_RAM_21 = 256'h7983D3C7C742032010B0FFBB8B175C8AFCE3F02EA0FA0000017206720175C012;
defparam prom_inst_1.INIT_RAM_22 = 256'hFBF572743C3C3C72743C727286FCE932F02E8E48B84D4AFFC30401E902C64933;
defparam prom_inst_1.INIT_RAM_23 = 256'hE903E6E4E61610409FBB33600780F4CD4AB8EB70260000D1000070B8A0741FCF;
defparam prom_inst_1.INIT_RAM_24 = 256'hEBF902F3CF0877FF000072F9EB00A4E8732A15061E06635D031C3CADE6E407C4;
defparam prom_inst_1.INIT_RAM_25 = 256'h0905781CFCEF86560000C828EBB4FF50028A9F92E8C5B48468D8AEE8E1B4B403;
defparam prom_inst_1.INIT_RAM_26 = 256'hE3C005EBE0808A7424B01C743B80723B898B1F0000E0363600AD8B16F4249212;
defparam prom_inst_1.INIT_RAM_27 = 256'hF724E812FA018EE7E64301F9BEEC08ECE000C8BAF780DB07E872E8F397720080;
defparam prom_inst_1.INIT_RAM_28 = 256'h00006E6C74FC6A00EACD0780B9002E303020623520536F69776C692076742000;
defparam prom_inst_1.INIT_RAM_29 = 256'hF9505006FC0067B368A4778B00D8006ACFE75B00530600839C74066AF98989FB;
defparam prom_inst_1.INIT_RAM_2A = 256'hFAFF72DBE4F108ECA8B7C3C4D4DBF108ECA8B7524242E9DCC0E80272EC03B407;
defparam prom_inst_1.INIT_RAM_2B = 256'hDAFFD1FFFFE99090EEB010C00EC30EFF74CAD200AFF52EEB9F001EAFCFAE10F6;
defparam prom_inst_1.INIT_RAM_2C = 256'hB5FCE8D8DEC1060AFF05168B01BA42F950F5EBC3FC46F6E8FF5BE225E8C3E201;
defparam prom_inst_1.INIT_RAM_2D = 256'hFEB5FC01B0D8DFC1060A8BFF051601BA42F950C38BEFF7E8D01FBEFD4BFF52D6;
defparam prom_inst_1.INIT_RAM_2E = 256'hCCE8FEA8F77558E88BB1FEF775D3F701FE0ABA51E9D0FEB88983F9FE750ED2E8;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000007A000069000049000040C15FEF8BC1FE162B75FE757CF774581FE1FEF1;
defparam prom_inst_1.INIT_RAM_30 = 256'h002F3F00003F3F001F3F3F382D28241C18140E0B08003F3F153F15152A2A002A;
defparam prom_inst_1.INIT_RAM_31 = 256'h15152A2A002A00002A2A002A00000E0A06021F3F3F1F2F3F10003F3F00003F1F;
defparam prom_inst_1.INIT_RAM_32 = 256'h153F15153F3F153F15152A2A002A00002A2A002A00003F3F153F15153F3F153F;
defparam prom_inst_1.INIT_RAM_33 = 256'h15003F2A153F00153F2A003F00002A2A152A00152A2A002A0000161206023F3F;
defparam prom_inst_1.INIT_RAM_34 = 256'h1509483C36313E3A14023F3F153F15153F3F003F15002A3F152A15152A3F002A;
defparam prom_inst_1.INIT_RAM_35 = 256'h1E1E1F1F2C2C10100000514C4548521C001E5456592C2E000013060019110443;
defparam prom_inst_1.INIT_RAM_36 = 256'h24243232151522222323303031311313141421212F2F121220202D2D2E2E1111;
defparam prom_inst_1.INIT_RAM_37 = 256'h844976518D48744D9150935392527747734B754F191926261818171725251616;
defparam prom_inst_1.INIT_RAM_38 = 256'h00040005030300020029940F613E6340654267448A865F3C5E3B603D623F8F4C;
defparam prom_inst_1.INIT_RAM_39 = 256'h000D1A1A00280C0C002795E000350034000A000B003300090008070700063939;
defparam prom_inst_1.INIT_RAM_3A = 256'h904E898501018D48744D66439150935392527747734B754F0E0E2B2B1B1B1C1C;
defparam prom_inst_1.INIT_RAM_3B = 256'h000000000000000000000000000000000000000064414646844996378E4A7651;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'hFF32315B00000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hE8E6F6E6E7E600BC300A74654B50642042657275616931295320434B6E673678;
defparam prom_inst_2.INIT_RAM_01 = 256'h48C7500AC748F8C7404AC720D4C7F608FE8CC7F61F75043CC0BAA5B933686815;
defparam prom_inst_2.INIT_RAM_02 = 256'h646410B884000984820003C744444413107803ABC0FF1FBEC7C064C764CBC758;
defparam prom_inst_2.INIT_RAM_03 = 256'hE4B0FB80B03C07F8E81913B486A8AD96730113B43C151372F2AA13E331E8FBE8;
defparam prom_inst_2.INIT_RAM_04 = 256'h65206F531603CD137104F6E07406E813D11386E807A3F8ECD2FB012100E6E68A;
defparam prom_inst_2.INIT_RAM_05 = 256'h0803C075C7C0803C07C51E2048692032444D4D0D62627A335031682030550D64;
defparam prom_inst_2.INIT_RAM_06 = 256'h4FE940EB00807514F63C8B8B406058EB747574E4FB0400000D3F1800016C6A58;
defparam prom_inst_2.INIT_RAM_07 = 256'h80C1B802378008F63CE2B60175EB0563803CC10034C70380E2530175EB050172;
defparam prom_inst_2.INIT_RAM_08 = 256'hC202A61BA300003EF67421FF100140FE628008F63C04EB0474130174193381E2;
defparam prom_inst_2.INIT_RAM_09 = 256'hB3C202F6022077EB13F63C74DBFA223CC1800B76F200FA85807422BF20E806F6;
defparam prom_inst_2.INIT_RAM_0A = 256'h078BFC4F40FC3280D4F309CF00000FB3327510C5C0E180055119001677FA2EE0;
defparam prom_inst_2.INIT_RAM_0B = 256'hEB0AFB1E808ACD8ACDFF7502EB2EBE5701F94F59C0A50ABEEB4F030D77CFBE01;
defparam prom_inst_2.INIT_RAM_0C = 256'hC487870202E6A00000016874446C4E00000000565883CBEF080A83018B9C0EDC;
defparam prom_inst_2.INIT_RAM_0D = 256'h00068FC7C73CC7C74C28C7141AE96914BEB800C74A0642432E58FF05B0B8080F;
defparam prom_inst_2.INIT_RAM_0E = 256'h49F6B9F706000006DFC74AF706BF4C28C775EB0402BA000006DF757420002200;
defparam prom_inst_2.INIT_RAM_0F = 256'h0606B4231100B02EEEC00375CD7559FF8E0059000050EFEF07B0EF8B07DCB824;
defparam prom_inst_2.INIT_RAM_10 = 256'h07C3EFEF8ABAC0C0753A0050E3C150EFEFB0C50485605010BBCD81CD69401075;
defparam prom_inst_2.INIT_RAM_11 = 256'h843ED200E8CAC3E7B0D4A3D8084C0A12E70A04CDCDE700777349A22460C30E8B;
defparam prom_inst_2.INIT_RAM_12 = 256'h07E8535803C7D88BB807508B53F0D1FA6B33EBF741F7C379038AE3CCF2F3032A;
defparam prom_inst_2.INIT_RAM_13 = 256'hB853763AB2B2D280594A10B93C3C3C3C00065B02E8E38BB78AC3E207E8E35BAB;
defparam prom_inst_2.INIT_RAM_14 = 256'hF260C78AEC60940377917258401069696969CFBA698E6900000080A05A331636;
defparam prom_inst_2.INIT_RAM_15 = 256'hC3C18A42BA52B70010AACDB3C38A42030352892432E6EE24E3A0B0EC6079108A;
defparam prom_inst_2.INIT_RAM_16 = 256'h3AC30352EE936C6B93FA58C88AEC038A61EEE7C058502ED0752EC0DA6103EEBA;
defparam prom_inst_2.INIT_RAM_17 = 256'hBABA0110E60000F7B86AA84B26F5BACBC3CF10CED11CB569F2C1B02BEF07E71E;
defparam prom_inst_2.INIT_RAM_18 = 256'h0EB8723EB884ACF6E3448933100733EC2E60D908C33C3C3C7274747474582E10;
defparam prom_inst_2.INIT_RAM_19 = 256'h243275C30F8875C8BAD8C3D3F6C177C3C47C0001848561DC10C87400006084F7;
defparam prom_inst_2.INIT_RAM_1A = 256'hBB0001B70210BBB82180ABEDC389BB8A3CCD74445850004546A85003F3E3C389;
defparam prom_inst_2.INIT_RAM_1B = 256'h0040253E252525E35C9B258A4EE78B46700001200C6133022400AB893300753E;
defparam prom_inst_2.INIT_RAM_1C = 256'hEFEFEFEFEFEEEFEFEEEEEE5D46D0F63626551E81E8AA0122EC1AFB001F1E136A;
defparam prom_inst_2.INIT_RAM_1D = 256'hC02B51E860C14A808403BD3274006A80FF8D921F06B4859475EFEFEFEFEFEFEE;
defparam prom_inst_2.INIT_RAM_1E = 256'h508037F6EBC3013FC0FE03F1B91EEAC194CB80AA80743ED2E2BA3FD2C1E1C3D8;
defparam prom_inst_2.INIT_RAM_1F = 256'hF26AC30000166C890A106C0C6C086C040B00ED8E9475C38061025E1E085C8B36;
defparam prom_inst_2.INIT_RAM_20 = 256'h40EDEB83A8EB8AFBECC3ECECEE4AC5EEEEE8B817C0EC8A525E5174088B7F8B14;
defparam prom_inst_2.INIT_RAM_21 = 256'h05DBFFF7778BC9071FFF4A04748B14648A72BA87F02E06A6EF033D0B830B8375;
defparam prom_inst_2.INIT_RAM_22 = 256'hCAB80362C09290E258862227C44F5EE46187164A02FF85E8748BA4F3A40174C0;
defparam prom_inst_2.INIT_RAM_23 = 256'h7D9DA1A164B8001F1ED6C07BEB7426150700C3F9A0B48900038C89E70021801E;
defparam prom_inst_2.INIT_RAM_24 = 256'hC5E858F9F22E8806EB8893E8A100C62CB0C7B8A3A174743C727401E6A1A177B4;
defparam prom_inst_2.INIT_RAM_25 = 256'h7474743CA874C46A0000083CAAE502EB72C8028AA602E9FF00128AC202F2E877;
defparam prom_inst_2.INIT_RAM_26 = 256'h1FE77597A0E4260277A000B7360004360C36CAAD3B8B1A80723B3674B45E7574;
defparam prom_inst_2.INIT_RAM_27 = 256'hEA460D018AE8C00142B8B00103C32A327424FADA5A26E88A110E99530023E8E3;
defparam prom_inst_2.INIT_RAM_28 = 256'h00C60000160140CD0013BB0001B82E293A66703228326E6E61656C61692062F0;
defparam prom_inst_2.INIT_RAM_29 = 256'h8353ACB474AD000000000CF0A0FEE440FC705080C5A0731E001BA040EB0E16CA;
defparam prom_inst_2.INIT_RAM_2A = 256'h757209E860C32A320128BAE6E674EB2A320228BA75385B73E808E8FAC0B9801F;
defparam prom_inst_2.INIT_RAM_2B = 256'hFF88E9E2ACACED9090FFEB74260ACD9203F52E00F52E8B400020B1F52EE67406;
defparam prom_inst_2.INIT_RAM_2C = 256'h02FEAC8303E81FE483FF1FD9EFDA5201B2500368FF74E8C4B9C3F60AC953F083;
defparam prom_inst_2.INIT_RAM_2D = 256'hE802E874FE8303E81FE4F383FF1FEFDA5201B250C5E85835ECE8DF01759DFF56;
defparam prom_inst_2.INIT_RAM_2E = 256'h74A2BEFE0E548091FC04CCE870FE0EEFE200DA5277ECE8FEB0FD4BD09880FED5;
defparam prom_inst_2.INIT_RAM_2F = 256'h2A00FF0000FF4000FF00019500595EE8E7C18B1FE114801CFE0E28A8E88BB1F7;
defparam prom_inst_2.INIT_RAM_30 = 256'h2F001F3F10003F3F00103F38322824201814110B08053F3F3F3F3F152A152A2A;
defparam prom_inst_2.INIT_RAM_31 = 256'h3F152A152A2A2A002A152A2A2A000F0B0703271F3F3F1F273F1F002F3F00003F;
defparam prom_inst_2.INIT_RAM_32 = 256'h3F3F3F153F3F3F3F3F152A152A2A2A002A152A2A2A003F3F3F3F3F153F3F3F3F;
defparam prom_inst_2.INIT_RAM_33 = 256'h2A153F3F2A3F3F002A3F2A2A3F003F2A2A3F2A002A2A2A2A2A00171307033F3F;
defparam prom_inst_2.INIT_RAM_34 = 256'h170D2F3B37323F3B07033F3F3F3F3F152A3F3F2A3F153F2A3F3F2A152A2A3F2A;
defparam prom_inst_2.INIT_RAM_35 = 256'h00410053005A00510000554D4951534F531F1B1C1D4F2628573A0A4740100346;
defparam prom_inst_2.INIT_RAM_36 = 256'h004A004D0059004700480042004E005200540046005600450044005800430057;
defparam prom_inst_2.INIT_RAM_37 = 256'h0A390433093807360332002E01300837053402310050004C004F0049004B0055;
defparam prom_inst_2.INIT_RAM_38 = 256'h0023002400400021007E00000000000000000000000000000000000000000635;
defparam prom_inst_2.INIT_RAM_39 = 256'h002B007B0022005F003A002F003F003E00280029003C002A0026005E00252020;
defparam prom_inst_2.INIT_RAM_3A = 256'h002B0000001B0000000000000000000000000000000000000008007C007D000D;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000002A002D0000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'hFF2F35E000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0DA1D04007439D0000FA657442530D43202B616D65633720204220206F2D2074;
defparam prom_inst_3.INIT_RAM_01 = 256'hF10600EE0600ED0600E30600E20689F3004C04BF1EF3060CEF80E800F6000000;
defparam prom_inst_3.INIT_RAM_02 = 256'hB9B0B0039671C787001E8344601C1A802403C7C7B1331EF40601F40600F30600;
defparam prom_inst_3.INIT_RAM_03 = 256'h6020E826A700E83C754972FF13E6E60005E872F083E83C1CE875722CB1E3B4D1;
defparam prom_inst_3.INIT_RAM_04 = 256'h63647532CD3314B8E27406E8069683BEE8A1E297BE94E8B4CDB440E6E76064E0;
defparam prom_inst_3.INIT_RAM_05 = 256'h5DC3E80200223FD8435E55004474314D52423A0A7569203653387A31313A0A0D;
defparam prom_inst_3.INIT_RAM_06 = 256'hF9AF8003E8E40CF6C5FA0E161F1E5B0204F60E64500100C7C7B07583830040CF;
defparam prom_inst_3.INIT_RAM_07 = 256'hE10275EB81CA80C138FE75EB055A803CCA2A02FF1206E9FC8075EB05EA803C03;
defparam prom_inst_3.INIT_RAM_08 = 256'h037500331CA380C6C745F60046733AEB81E280C19D01798008F63C1200C0E2F7;
defparam prom_inst_3.INIT_RAM_09 = 256'h0608B3C280750A0E80C21A02F62EC4590275EB26AEFC5100CE05F60045C6BBC2;
defparam prom_inst_3.INIT_RAM_0A = 256'h81F01C741F1EF3F9C3328A3207898900E80BF624E8FCE6CD8B00D58A0E838B03;
defparam prom_inst_3.INIT_RAM_0B = 256'hB3DF2549E73E10C310230A3DDDA55DB97501EBB4F3B10032E8B872743C3CED2E;
defparam prom_inst_3.INIT_RAM_0C = 256'h030000C00000004007FF6572756169F000F0014558E0ED5AE884E004C3FA6800;
defparam prom_inst_3.INIT_RAM_0D = 256'hC74AB4F8061CF8060000068F75AE008F20B910060008E6B0B03CEFEF0301EFEF;
defparam prom_inst_3.INIT_RAM_0E = 256'h00D000BB6900C74AB40074EB6928000006193B00FFC400C74AB420E3BF97C700;
defparam prom_inst_3.INIT_RAM_0F = 256'h89CD0111CDEE13A28A03ECEC10088051C380F605F30033B8121397C7BAFF090B;
defparam prom_inst_3.INIT_RAM_10 = 256'h83535A58E0D45086180603800EEB535A400ABA03000052070110C2100000331F;
defparam prom_inst_3.INIT_RAM_11 = 256'hDB4E03B8472B60480D034EC1F700E7758A00EB10108BE72519006207E8B46057;
defparam prom_inst_3.INIT_RAM_12 = 256'h87D951C3D86B335FC18D8107E8A08AB2F8C0B9DAE8D9FDF6FACB93790326F7E3;
defparam prom_inst_3.INIT_RAM_13 = 256'h0152E636000000EAC30042010D0A0807751858CD080757001E50F983C50E0787;
defparam prom_inst_3.INIT_RAM_14 = 256'hB3B0EEC3BABA24F609EBEBEBEBEBEAEAEAEAEAEAEAEAEAC38A8A0A875BC94A84;
defparam prom_inst_3.INIT_RAM_15 = 256'h60EEC58AC89200AA7543100060F8EC8AEC50002006C02EF7036F10BABAF54E7C;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFB3EC9393BA61C9EEBAC35AE88AEEC3C38A0272EBB0A2CF11A00303C3F342C8;
defparam prom_inst_3.INIT_RAM_17 = 256'hC0DA7532322E8848904010756EEFCBC16075FEB08A0300D24DEA156002750F6F;
defparam prom_inst_3.INIT_RAM_18 = 256'h85E01049C80E0C8EAB7E6CF60724D2B98BBBEC2E60302421EB1E1726AFC3A2EE;
defparam prom_inst_3.INIT_RAM_19 = 256'h08060F80BB000B80000000EC2EEE0E802E001F770000C3CD48B003D80E0600F1;
defparam prom_inst_3.INIT_RAM_1A = 256'h0113800003720808003CBEAB601E08C401100450E2E845260002B4F6C131B000;
defparam prom_inst_3.INIT_RAM_1B = 256'h1F1FE8EDE8E8E8ECEAE9E8E9E9E8E8E8E6000100608AC0AA07C0AB00C0AB0349;
defparam prom_inst_3.INIT_RAM_1C = 256'h9B2525F425D6252525D6CC1F085EDC9274EE2EE5C1EBEB762676FC0880550040;
defparam prom_inst_3.INIT_RAM_1D = 256'hD4C8FF12B43FB4FAC0BDB2F600C3EBFAB986001FC1FDC900298025F470BBC9F4;
defparam prom_inst_3.INIT_RAM_1E = 256'h6075F6EB08BDFE8BE0037648C18306E000B3B4C37405940003C1033FEAC08A61;
defparam prom_inst_3.INIT_RAM_1F = 256'h03401EC302C71444C1C10E3F0AFF06FF00C7C75E008580E458011F568B044C8E;
defparam prom_inst_3.INIT_RAM_20 = 256'h8325F1C201E8C483A852864A594A244242830004E90CE8515A4E4374C6EEF083;
defparam prom_inst_3.INIT_RAM_21 = 256'h03002BD802C61333686893E8127C8A1F440682260E8C1EF0C32D0083F825F802;
defparam prom_inst_3.INIT_RAM_22 = 256'h0200743C727272743C72743C3C74FFEB1F26A0EF00EBF6530DC8E8A549000F43;
defparam prom_inst_3.INIT_RAM_23 = 256'hFF5AE824F9A704F652F20EEBAAF9F672338306F500010EA3C2061E037584F46A;
defparam prom_inst_3.INIT_RAM_24 = 256'h80F372E8508AC1B4E63EBB1BB43206038A38F500007527054033FA64FB0CE701;
defparam prom_inst_3.INIT_RAM_25 = 256'h083D7B03EF3E4840001000500A02778284E872D80272F975EBC7F80272F9EBDF;
defparam prom_inst_3.INIT_RAM_26 = 256'h0A059280170C962CA81848891AB08B82461C02FB3636000004361AF9111F0256;
defparam prom_inst_3.INIT_RAM_27 = 256'h004B018AFC18BE8EE600B4E8F40EF8C70A58A003EB9788E300B401320880287F;
defparam prom_inst_3.INIT_RAM_28 = 256'hF506A08B8B771F187C72006A00010D203130733031332067692C617663646F4E;
defparam prom_inst_3.INIT_RAM_29 = 256'hC4FF5000120BBE88753A882C6706601F6058330F1E00149EE881001FEA6E6C02;
defparam prom_inst_3.INIT_RAM_2A = 256'hF704E8BCC3A8F8C775E4DA6064040CF8C774E4DAF8E80AF50200E4E4E852BA61;
defparam prom_inst_3.INIT_RAM_2B = 256'h8825E8F6E8E8C39090B4F404AC001005E885F75200FF1E75BF2EF52E8F640496;
defparam prom_inst_3.INIT_RAM_2C = 256'h5E75FFE7C6048B75C4E8C68B8B038B74518A680A7405B0FF06E8F6DCFF320BC7;
defparam prom_inst_3.INIT_RAM_2D = 256'hD8E8E20283E6C7048B758BC4E8C68B038B74588A2B2C33FF7381F774D772E89C;
defparam prom_inst_3.INIT_RAM_2E = 256'hEBFEE5E81FBEFCFE162B75C6BEFE1FBEFBE80356FF73B0E8FD0175ECE8FC80FE;
defparam prom_inst_3.INIT_RAM_2F = 256'h00000000007700004C00AA48001F5A1433084DE88BB1FCE80A1FBE4064FC04E8;
defparam prom_inst_3.INIT_RAM_30 = 256'h3F3F00103F1F003F3F000038322D24201C14110E08050015153F15151500002A;
defparam prom_inst_3.INIT_RAM_31 = 256'h15151500002A00000000002A0000000C0804002F1F3F3F1F1F3F2F001F3F0000;
defparam prom_inst_3.INIT_RAM_32 = 256'h153F15151515153F15151500002A00000000002A00000015153F15151515153F;
defparam prom_inst_3.INIT_RAM_33 = 256'h00001515152A15150000152A00150015002A15000000002A0000001410040015;
defparam prom_inst_3.INIT_RAM_34 = 256'h180C01413834003C38040015153F15151500153F00151515003F15001500003F;
defparam prom_inst_3.INIT_RAM_35 = 256'h1E1E1F1F2C2C10100000584E4A49504B2A002025222B2D29003D0F0242140845;
defparam prom_inst_3.INIT_RAM_36 = 256'h24243232151522222323303031311313141421212F2F121220202D2D2E2E1111;
defparam prom_inst_3.INIT_RAM_37 = 256'h004900510048004D0050005300520047004B004F191926261818171725251616;
defparam prom_inst_3.INIT_RAM_38 = 256'h7A047B05790378022929000F6B576D596F5B715D8C88695568546A566C58004C;
defparam prom_inst_3.INIT_RAM_39 = 256'h830D1A1A2828820C2727A4E035353434800A810B33337F097E087D077C063939;
defparam prom_inst_3.INIT_RAM_3A = 256'h4E4E8B87010198489D4D705CA050A353A25297479B4B9F4F0E0E2B2B1B1B1C1C;
defparam prom_inst_3.INIT_RAM_3B = 256'h00000000000000000000000000000000000000006E5A4646994937374A4AA151;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h00312F0000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_pROM_bios
