//-----------------------------------------------------------------------------
//
// RAM image for input code file: hello.hex
//
//-----------------------------------------------------------------------------
module ram_image
(
	clk, addr, 
	we, din, dout
);
//-----------------------------------------------------------------------------
input           clk;
input   [12:0]  addr;
input           we;
input   [7:0]   din;
output  [7:0]   dout;
//-----------------------------------------------------------------------------
reg [7:0] dout;
reg [7:0] ram [8191:0];
//-----------------------------------------------------------------------------
initial 
begin
	ram[0] = 8'hf3;	ram[1] = 8'hc3;	ram[2] = 8'h21;	ram[3] = 8'h0d;
	ram[4] = 8'h90;	ram[5] = 8'h04;	ram[6] = 8'hf9;	ram[7] = 8'h07;
	ram[8] = 8'h7e;	ram[9] = 8'he3;	ram[10] = 8'hbe;	ram[11] = 8'h23;
	ram[12] = 8'he3;	ram[13] = 8'hc2;	ram[14] = 8'hd0;	ram[15] = 8'h01;
	ram[16] = 8'h23;	ram[17] = 8'h7e;	ram[18] = 8'hfe;	ram[19] = 8'h3a;
	ram[20] = 8'hd0;	ram[21] = 8'hc3;	ram[22] = 8'h5e;	ram[23] = 8'h04;
	ram[24] = 8'hf5;	ram[25] = 8'h3a;	ram[26] = 8'h27;	ram[27] = 8'h00;
	ram[28] = 8'hc3;	ram[29] = 8'h6e;	ram[30] = 8'h03;	ram[31] = 8'h00;
	ram[32] = 8'h7c;	ram[33] = 8'h92;	ram[34] = 8'hc0;	ram[35] = 8'h7d;
	ram[36] = 8'h93;	ram[37] = 8'hc9;	ram[38] = 8'h01;	ram[39] = 8'h00;
	ram[40] = 8'h3a;	ram[41] = 8'h72;	ram[42] = 8'h01;	ram[43] = 8'hb7;
	ram[44] = 8'hc2;	ram[45] = 8'hda;	ram[46] = 8'h09;	ram[47] = 8'hc9;
	ram[48] = 8'he3;	ram[49] = 8'h22;	ram[50] = 8'h3b;	ram[51] = 8'h00;
	ram[52] = 8'he1;	ram[53] = 8'h4e;	ram[54] = 8'h23;	ram[55] = 8'h46;
	ram[56] = 8'h23;	ram[57] = 8'hc5;	ram[58] = 8'hc3;	ram[59] = 8'h3a;
	ram[60] = 8'h00;	ram[61] = 8'he4;	ram[62] = 8'h09;	ram[63] = 8'ha2;
	ram[64] = 8'h0a;	ram[65] = 8'hf8;	ram[66] = 8'h09;	ram[67] = 8'h98;
	ram[68] = 8'h04;	ram[69] = 8'h21;	ram[70] = 8'h0c;	ram[71] = 8'h5f;
	ram[72] = 8'h0c;	ram[73] = 8'h95;	ram[74] = 8'h0c;	ram[75] = 8'h79;
	ram[76] = 8'h10;	ram[77] = 8'h08;	ram[78] = 8'h79;	ram[79] = 8'h0a;
	ram[80] = 8'h08;	ram[81] = 8'h7c;	ram[82] = 8'he3;	ram[83] = 8'h08;
	ram[84] = 8'h7c;	ram[85] = 8'h2f;	ram[86] = 8'h09;	ram[87] = 8'h45;
	ram[88] = 8'h4e;	ram[89] = 8'hc4;	ram[90] = 8'h46;	ram[91] = 8'h4f;
	ram[92] = 8'hd2;	ram[93] = 8'h4e;	ram[94] = 8'h45;	ram[95] = 8'h58;
	ram[96] = 8'hd4;	ram[97] = 8'h44;	ram[98] = 8'h41;	ram[99] = 8'h54;
	ram[100] = 8'hc1;	ram[101] = 8'h49;	ram[102] = 8'h4e;	ram[103] = 8'h50;
	ram[104] = 8'h55;	ram[105] = 8'hd4;	ram[106] = 8'h44;	ram[107] = 8'h49;
	ram[108] = 8'hcd;	ram[109] = 8'h52;	ram[110] = 8'h45;	ram[111] = 8'h41;
	ram[112] = 8'hc4;	ram[113] = 8'h4c;	ram[114] = 8'h45;	ram[115] = 8'hd4;
	ram[116] = 8'h47;	ram[117] = 8'h4f;	ram[118] = 8'h54;	ram[119] = 8'hcf;
	ram[120] = 8'h52;	ram[121] = 8'h55;	ram[122] = 8'hce;	ram[123] = 8'h49;
	ram[124] = 8'hc6;	ram[125] = 8'h52;	ram[126] = 8'h45;	ram[127] = 8'h53;
	ram[128] = 8'h54;	ram[129] = 8'h4f;	ram[130] = 8'h52;	ram[131] = 8'hc5;
	ram[132] = 8'h47;	ram[133] = 8'h4f;	ram[134] = 8'h53;	ram[135] = 8'h55;
	ram[136] = 8'hc2;	ram[137] = 8'h52;	ram[138] = 8'h45;	ram[139] = 8'h54;
	ram[140] = 8'h55;	ram[141] = 8'h52;	ram[142] = 8'hce;	ram[143] = 8'h52;
	ram[144] = 8'h45;	ram[145] = 8'hcd;	ram[146] = 8'h53;	ram[147] = 8'h54;
	ram[148] = 8'h4f;	ram[149] = 8'hd0;	ram[150] = 8'h50;	ram[151] = 8'h52;
	ram[152] = 8'h49;	ram[153] = 8'h4e;	ram[154] = 8'hd4;	ram[155] = 8'h4c;
	ram[156] = 8'h49;	ram[157] = 8'h53;	ram[158] = 8'hd4;	ram[159] = 8'h43;
	ram[160] = 8'h4c;	ram[161] = 8'h45;	ram[162] = 8'h41;	ram[163] = 8'hd2;
	ram[164] = 8'h4e;	ram[165] = 8'h45;	ram[166] = 8'hd7;	ram[167] = 8'h54;
	ram[168] = 8'h41;	ram[169] = 8'h42;	ram[170] = 8'ha8;	ram[171] = 8'h54;
	ram[172] = 8'hcf;	ram[173] = 8'h54;	ram[174] = 8'h48;	ram[175] = 8'h45;
	ram[176] = 8'hce;	ram[177] = 8'h53;	ram[178] = 8'h54;	ram[179] = 8'h45;
	ram[180] = 8'hd0;	ram[181] = 8'hab;	ram[182] = 8'had;	ram[183] = 8'haa;
	ram[184] = 8'haf;	ram[185] = 8'hbe;	ram[186] = 8'hbd;	ram[187] = 8'hbc;
	ram[188] = 8'h53;	ram[189] = 8'h47;	ram[190] = 8'hce;	ram[191] = 8'h49;
	ram[192] = 8'h4e;	ram[193] = 8'hd4;	ram[194] = 8'h41;	ram[195] = 8'h42;
	ram[196] = 8'hd3;	ram[197] = 8'h55;	ram[198] = 8'h53;	ram[199] = 8'hd2;
	ram[200] = 8'h53;	ram[201] = 8'h51;	ram[202] = 8'hd2;	ram[203] = 8'h52;
	ram[204] = 8'h4e;	ram[205] = 8'hc4;	ram[206] = 8'h53;	ram[207] = 8'h49;
	ram[208] = 8'hce;	ram[209] = 8'h00;	ram[210] = 8'hf7;	ram[211] = 8'h01;
	ram[212] = 8'hd5;	ram[213] = 8'h03;	ram[214] = 8'h49;	ram[215] = 8'h06;
	ram[216] = 8'hf5;	ram[217] = 8'h04;	ram[218] = 8'he4;	ram[219] = 8'h05;
	ram[220] = 8'h16;	ram[221] = 8'h07;	ram[222] = 8'hf6;	ram[223] = 8'h05;
	ram[224] = 8'h02;	ram[225] = 8'h05;	ram[226] = 8'hcf;	ram[227] = 8'h04;
	ram[228] = 8'ha1;	ram[229] = 8'h02;	ram[230] = 8'h16;	ram[231] = 8'h05;
	ram[232] = 8'h69;	ram[233] = 8'h04;	ram[234] = 8'hbe;	ram[235] = 8'h04;
	ram[236] = 8'hdf;	ram[237] = 8'h04;	ram[238] = 8'hf7;	ram[239] = 8'h04;
	ram[240] = 8'hf7;	ram[241] = 8'h01;	ram[242] = 8'h57;	ram[243] = 8'h05;
	ram[244] = 8'h8e;	ram[245] = 8'h03;	ram[246] = 8'ha6;	ram[247] = 8'h02;
	ram[248] = 8'h95;	ram[249] = 8'h02;	ram[250] = 8'h4e;	ram[251] = 8'hc6;
	ram[252] = 8'h53;	ram[253] = 8'hce;	ram[254] = 8'h52;	ram[255] = 8'hc7;
	ram[256] = 8'h4f;	ram[257] = 8'hc4;	ram[258] = 8'h46;	ram[259] = 8'hc3;
	ram[260] = 8'h4f;	ram[261] = 8'hd6;	ram[262] = 8'h4f;	ram[263] = 8'hcd;
	ram[264] = 8'h55;	ram[265] = 8'hd3;	ram[266] = 8'h42;	ram[267] = 8'hd3;
	ram[268] = 8'h44;	ram[269] = 8'hc4;	ram[270] = 8'h2f;	ram[271] = 8'hb0;
	ram[272] = 8'h49;	ram[273] = 8'hc4;	ram[274] = 8'h2c;	ram[275] = 8'h00;
	ram[276] = 8'h00;	ram[277] = 8'h00;	ram[278] = 8'h00;	ram[279] = 8'h00;
	ram[280] = 8'h00;	ram[281] = 8'h00;	ram[282] = 8'h00;	ram[283] = 8'h00;
	ram[284] = 8'h00;	ram[285] = 8'h00;	ram[286] = 8'h00;	ram[287] = 8'h00;
	ram[288] = 8'h00;	ram[289] = 8'h00;	ram[290] = 8'h00;	ram[291] = 8'h00;
	ram[292] = 8'h00;	ram[293] = 8'h00;	ram[294] = 8'h00;	ram[295] = 8'h00;
	ram[296] = 8'h00;	ram[297] = 8'h00;	ram[298] = 8'h00;	ram[299] = 8'h00;
	ram[300] = 8'h00;	ram[301] = 8'h00;	ram[302] = 8'h00;	ram[303] = 8'h00;
	ram[304] = 8'h00;	ram[305] = 8'h00;	ram[306] = 8'h00;	ram[307] = 8'h00;
	ram[308] = 8'h00;	ram[309] = 8'h00;	ram[310] = 8'h00;	ram[311] = 8'h00;
	ram[312] = 8'h00;	ram[313] = 8'h00;	ram[314] = 8'h00;	ram[315] = 8'h00;
	ram[316] = 8'h00;	ram[317] = 8'h00;	ram[318] = 8'h00;	ram[319] = 8'h00;
	ram[320] = 8'h00;	ram[321] = 8'h00;	ram[322] = 8'h00;	ram[323] = 8'h00;
	ram[324] = 8'h00;	ram[325] = 8'h00;	ram[326] = 8'h00;	ram[327] = 8'h00;
	ram[328] = 8'h00;	ram[329] = 8'h00;	ram[330] = 8'h00;	ram[331] = 8'h00;
	ram[332] = 8'h00;	ram[333] = 8'h00;	ram[334] = 8'h00;	ram[335] = 8'h00;
	ram[336] = 8'h00;	ram[337] = 8'h00;	ram[338] = 8'h00;	ram[339] = 8'h00;
	ram[340] = 8'h00;	ram[341] = 8'h00;	ram[342] = 8'h00;	ram[343] = 8'h00;
	ram[344] = 8'h00;	ram[345] = 8'h00;	ram[346] = 8'h00;	ram[347] = 8'h00;
	ram[348] = 8'h00;	ram[349] = 8'h00;	ram[350] = 8'h00;	ram[351] = 8'h00;
	ram[352] = 8'h00;	ram[353] = 8'h00;	ram[354] = 8'h00;	ram[355] = 8'h1a;
	ram[356] = 8'h0f;	ram[357] = 8'h00;	ram[358] = 8'h00;	ram[359] = 8'h00;
	ram[360] = 8'h00;	ram[361] = 8'h00;	ram[362] = 8'h00;	ram[363] = 8'h00;
	ram[364] = 8'h00;	ram[365] = 8'h00;	ram[366] = 8'h00;	ram[367] = 8'h00;
	ram[368] = 8'h00;	ram[369] = 8'h00;	ram[370] = 8'h00;	ram[371] = 8'h00;
	ram[372] = 8'h00;	ram[373] = 8'h00;	ram[374] = 8'h00;	ram[375] = 8'h00;
	ram[376] = 8'h00;	ram[377] = 8'h00;	ram[378] = 8'h00;	ram[379] = 8'h00;
	ram[380] = 8'h00;	ram[381] = 8'h00;	ram[382] = 8'h00;	ram[383] = 8'h00;
	ram[384] = 8'h00;	ram[385] = 8'h20;	ram[386] = 8'h45;	ram[387] = 8'h52;
	ram[388] = 8'h52;	ram[389] = 8'h4f;	ram[390] = 8'hd2;	ram[391] = 8'h00;
	ram[392] = 8'h20;	ram[393] = 8'h49;	ram[394] = 8'h4e;	ram[395] = 8'ha0;
	ram[396] = 8'h00;	ram[397] = 8'h0d;	ram[398] = 8'h4f;	ram[399] = 8'hcb;
	ram[400] = 8'h0d;	ram[401] = 8'h00;	ram[402] = 8'h21;	ram[403] = 8'h04;
	ram[404] = 8'h00;	ram[405] = 8'h39;	ram[406] = 8'h7e;	ram[407] = 8'h23;
	ram[408] = 8'hfe;	ram[409] = 8'h81;	ram[410] = 8'hc0;	ram[411] = 8'hf7;
	ram[412] = 8'he3;	ram[413] = 8'he7;	ram[414] = 8'h01;	ram[415] = 8'h0d;
	ram[416] = 8'h00;	ram[417] = 8'he1;	ram[418] = 8'hc8;	ram[419] = 8'h09;
	ram[420] = 8'hc3;	ram[421] = 8'h96;	ram[422] = 8'h01;	ram[423] = 8'hcd;
	ram[424] = 8'hc3;	ram[425] = 8'h01;	ram[426] = 8'hc5;	ram[427] = 8'he3;
	ram[428] = 8'hc1;	ram[429] = 8'he7;	ram[430] = 8'h7e;	ram[431] = 8'h02;
	ram[432] = 8'hc8;	ram[433] = 8'h0b;	ram[434] = 8'h2b;	ram[435] = 8'hc3;
	ram[436] = 8'had;	ram[437] = 8'h01;	ram[438] = 8'he5;	ram[439] = 8'h2a;
	ram[440] = 8'h6b;	ram[441] = 8'h01;	ram[442] = 8'h06;	ram[443] = 8'h00;
	ram[444] = 8'h09;	ram[445] = 8'h09;	ram[446] = 8'hcd;	ram[447] = 8'hc3;
	ram[448] = 8'h01;	ram[449] = 8'he1;	ram[450] = 8'hc9;	ram[451] = 8'hd5;
	ram[452] = 8'heb;	ram[453] = 8'h21;	ram[454] = 8'hde;	ram[455] = 8'hff;
	ram[456] = 8'h39;	ram[457] = 8'he7;	ram[458] = 8'heb;	ram[459] = 8'hd1;
	ram[460] = 8'hd0;	ram[461] = 8'h1e;	ram[462] = 8'h0c;	ram[463] = 8'h01;
	ram[464] = 8'h1e;	ram[465] = 8'h02;	ram[466] = 8'h01;	ram[467] = 8'h1e;
	ram[468] = 8'h14;	ram[469] = 8'hcd;	ram[470] = 8'hb5;	ram[471] = 8'h02;
	ram[472] = 8'hcd;	ram[473] = 8'h8a;	ram[474] = 8'h05;	ram[475] = 8'h21;
	ram[476] = 8'hfa;	ram[477] = 8'h00;	ram[478] = 8'h57;	ram[479] = 8'h3e;
	ram[480] = 8'h3f;	ram[481] = 8'hdf;	ram[482] = 8'h19;	ram[483] = 8'h7e;
	ram[484] = 8'hdf;	ram[485] = 8'hd7;	ram[486] = 8'hdf;	ram[487] = 8'h21;
	ram[488] = 8'h81;	ram[489] = 8'h01;	ram[490] = 8'hcd;	ram[491] = 8'ha3;
	ram[492] = 8'h05;	ram[493] = 8'h2a;	ram[494] = 8'h61;	ram[495] = 8'h01;
	ram[496] = 8'h7c;	ram[497] = 8'ha5;	ram[498] = 8'h3c;	ram[499] = 8'hc4;
	ram[500] = 8'h2f;	ram[501] = 8'h0b;	ram[502] = 8'h01;	ram[503] = 8'hc0;
	ram[504] = 8'hc1;	ram[505] = 8'h21;	ram[506] = 8'h8d;	ram[507] = 8'h01;
	ram[508] = 8'hcd;	ram[509] = 8'h21;	ram[510] = 8'h0d;	ram[511] = 8'h21;
	ram[512] = 8'hff;	ram[513] = 8'hff;	ram[514] = 8'h22;	ram[515] = 8'h61;
	ram[516] = 8'h01;	ram[517] = 8'hcd;	ram[518] = 8'h3c;	ram[519] = 8'h03;
	ram[520] = 8'hd7;	ram[521] = 8'h3c;	ram[522] = 8'h3d;	ram[523] = 8'hca;
	ram[524] = 8'hff;	ram[525] = 8'h01;	ram[526] = 8'hf5;	ram[527] = 8'hcd;
	ram[528] = 8'h9d;	ram[529] = 8'h04;	ram[530] = 8'hd5;	ram[531] = 8'hcd;
	ram[532] = 8'hcc;	ram[533] = 8'h02;	ram[534] = 8'h47;	ram[535] = 8'hd1;
	ram[536] = 8'hf1;	ram[537] = 8'hd2;	ram[538] = 8'h3e;	ram[539] = 8'h04;
	ram[540] = 8'hd5;	ram[541] = 8'hc5;	ram[542] = 8'hd7;	ram[543] = 8'hb7;
	ram[544] = 8'hf5;	ram[545] = 8'hcd;	ram[546] = 8'h7d;	ram[547] = 8'h02;
	ram[548] = 8'hc5;	ram[549] = 8'hd2;	ram[550] = 8'h39;	ram[551] = 8'h02;
	ram[552] = 8'heb;	ram[553] = 8'h2a;	ram[554] = 8'h67;	ram[555] = 8'h01;
	ram[556] = 8'h1a;	ram[557] = 8'h02;	ram[558] = 8'h03;	ram[559] = 8'h13;
	ram[560] = 8'he7;	ram[561] = 8'hc2;	ram[562] = 8'h2c;	ram[563] = 8'h02;
	ram[564] = 8'h60;	ram[565] = 8'h69;	ram[566] = 8'h22;	ram[567] = 8'h67;
	ram[568] = 8'h01;	ram[569] = 8'hd1;	ram[570] = 8'hf1;	ram[571] = 8'hca;
	ram[572] = 8'h60;	ram[573] = 8'h02;	ram[574] = 8'h2a;	ram[575] = 8'h67;
	ram[576] = 8'h01;	ram[577] = 8'he3;	ram[578] = 8'hc1;	ram[579] = 8'h09;
	ram[580] = 8'he5;	ram[581] = 8'hcd;	ram[582] = 8'ha7;	ram[583] = 8'h01;
	ram[584] = 8'he1;	ram[585] = 8'h22;	ram[586] = 8'h67;	ram[587] = 8'h01;
	ram[588] = 8'heb;	ram[589] = 8'h74;	ram[590] = 8'h23;	ram[591] = 8'h23;
	ram[592] = 8'hd1;	ram[593] = 8'h73;	ram[594] = 8'h23;	ram[595] = 8'h72;
	ram[596] = 8'h23;	ram[597] = 8'h11;	ram[598] = 8'h13;	ram[599] = 8'h01;
	ram[600] = 8'h1a;	ram[601] = 8'h77;	ram[602] = 8'h23;	ram[603] = 8'h13;
	ram[604] = 8'hb7;	ram[605] = 8'hc2;	ram[606] = 8'h58;	ram[607] = 8'h02;
	ram[608] = 8'hcd;	ram[609] = 8'ha2;	ram[610] = 8'h02;	ram[611] = 8'h23;
	ram[612] = 8'heb;	ram[613] = 8'h62;	ram[614] = 8'h6b;	ram[615] = 8'h7e;
	ram[616] = 8'h23;	ram[617] = 8'hb6;	ram[618] = 8'hca;	ram[619] = 8'hff;
	ram[620] = 8'h01;	ram[621] = 8'h23;	ram[622] = 8'h23;	ram[623] = 8'h23;
	ram[624] = 8'haf;	ram[625] = 8'hbe;	ram[626] = 8'h23;	ram[627] = 8'hc2;
	ram[628] = 8'h71;	ram[629] = 8'h02;	ram[630] = 8'heb;	ram[631] = 8'h73;
	ram[632] = 8'h23;	ram[633] = 8'h72;	ram[634] = 8'hc3;	ram[635] = 8'h65;
	ram[636] = 8'h02;	ram[637] = 8'h2a;	ram[638] = 8'h65;	ram[639] = 8'h01;
	ram[640] = 8'h44;	ram[641] = 8'h4d;	ram[642] = 8'h7e;	ram[643] = 8'h23;
	ram[644] = 8'hb6;	ram[645] = 8'h2b;	ram[646] = 8'hc8;	ram[647] = 8'hc5;
	ram[648] = 8'hf7;	ram[649] = 8'hf7;	ram[650] = 8'he1;	ram[651] = 8'he7;
	ram[652] = 8'he1;	ram[653] = 8'hc1;	ram[654] = 8'h3f;	ram[655] = 8'hc8;
	ram[656] = 8'h3f;	ram[657] = 8'hd0;	ram[658] = 8'hc3;	ram[659] = 8'h80;
	ram[660] = 8'h02;	ram[661] = 8'hc0;	ram[662] = 8'h2a;	ram[663] = 8'h65;
	ram[664] = 8'h01;	ram[665] = 8'haf;	ram[666] = 8'h77;	ram[667] = 8'h23;
	ram[668] = 8'h77;	ram[669] = 8'h23;	ram[670] = 8'h22;	ram[671] = 8'h67;
	ram[672] = 8'h01;	ram[673] = 8'hc0;	ram[674] = 8'h2a;	ram[675] = 8'h65;
	ram[676] = 8'h01;	ram[677] = 8'h2b;	ram[678] = 8'h22;	ram[679] = 8'h5d;
	ram[680] = 8'h01;	ram[681] = 8'hcd;	ram[682] = 8'h69;	ram[683] = 8'h04;
	ram[684] = 8'h2a;	ram[685] = 8'h67;	ram[686] = 8'h01;	ram[687] = 8'h22;
	ram[688] = 8'h69;	ram[689] = 8'h01;	ram[690] = 8'h22;	ram[691] = 8'h6b;
	ram[692] = 8'h01;	ram[693] = 8'hc1;	ram[694] = 8'h2a;	ram[695] = 8'h63;
	ram[696] = 8'h01;	ram[697] = 8'hf9;	ram[698] = 8'haf;	ram[699] = 8'h6f;
	ram[700] = 8'he5;	ram[701] = 8'hc5;	ram[702] = 8'h2a;	ram[703] = 8'h5d;
	ram[704] = 8'h01;	ram[705] = 8'hc9;	ram[706] = 8'h3e;	ram[707] = 8'h3f;
	ram[708] = 8'hdf;	ram[709] = 8'h3e;	ram[710] = 8'h20;	ram[711] = 8'hdf;
	ram[712] = 8'hcd;	ram[713] = 8'h3c;	ram[714] = 8'h03;	ram[715] = 8'h23;
	ram[716] = 8'h0e;	ram[717] = 8'h05;	ram[718] = 8'h11;	ram[719] = 8'h13;
	ram[720] = 8'h01;	ram[721] = 8'h7e;	ram[722] = 8'hfe;	ram[723] = 8'h20;
	ram[724] = 8'hca;	ram[725] = 8'h02;	ram[726] = 8'h03;	ram[727] = 8'h47;
	ram[728] = 8'hfe;	ram[729] = 8'h22;	ram[730] = 8'hca;	ram[731] = 8'h15;
	ram[732] = 8'h03;	ram[733] = 8'hb7;	ram[734] = 8'hca;	ram[735] = 8'h29;
	ram[736] = 8'h03;	ram[737] = 8'hd5;	ram[738] = 8'h06;	ram[739] = 8'h00;
	ram[740] = 8'h11;	ram[741] = 8'h56;	ram[742] = 8'h00;	ram[743] = 8'he5;
	ram[744] = 8'h3e;	ram[745] = 8'hd7;	ram[746] = 8'h13;	ram[747] = 8'h1a;
	ram[748] = 8'he6;	ram[749] = 8'h7f;	ram[750] = 8'hca;	ram[751] = 8'hff;
	ram[752] = 8'h02;	ram[753] = 8'hbe;	ram[754] = 8'hc2;	ram[755] = 8'h1c;
	ram[756] = 8'h03;	ram[757] = 8'h1a;	ram[758] = 8'hb7;	ram[759] = 8'hf2;
	ram[760] = 8'he9;	ram[761] = 8'h02;	ram[762] = 8'hf1;	ram[763] = 8'h78;
	ram[764] = 8'hf6;	ram[765] = 8'h80;	ram[766] = 8'hf2;	ram[767] = 8'he1;
	ram[768] = 8'h7e;	ram[769] = 8'hd1;	ram[770] = 8'h23;	ram[771] = 8'h12;
	ram[772] = 8'h13;	ram[773] = 8'h0c;	ram[774] = 8'hd6;	ram[775] = 8'h8e;
	ram[776] = 8'hc2;	ram[777] = 8'hd1;	ram[778] = 8'h02;	ram[779] = 8'h47;
	ram[780] = 8'h7e;	ram[781] = 8'hb7;	ram[782] = 8'hca;	ram[783] = 8'h29;
	ram[784] = 8'h03;	ram[785] = 8'hb8;	ram[786] = 8'hca;	ram[787] = 8'h02;
	ram[788] = 8'h03;	ram[789] = 8'h23;	ram[790] = 8'h12;	ram[791] = 8'h0c;
	ram[792] = 8'h13;	ram[793] = 8'hc3;	ram[794] = 8'h0c;	ram[795] = 8'h03;
	ram[796] = 8'he1;	ram[797] = 8'he5;	ram[798] = 8'h04;	ram[799] = 8'heb;
	ram[800] = 8'hb6;	ram[801] = 8'h23;	ram[802] = 8'hf2;	ram[803] = 8'h20;
	ram[804] = 8'h03;	ram[805] = 8'heb;	ram[806] = 8'hc3;	ram[807] = 8'heb;
	ram[808] = 8'h02;	ram[809] = 8'h21;	ram[810] = 8'h12;	ram[811] = 8'h01;
	ram[812] = 8'h12;	ram[813] = 8'h13;	ram[814] = 8'h12;	ram[815] = 8'h13;
	ram[816] = 8'h12;	ram[817] = 8'hc9;	ram[818] = 8'h05;	ram[819] = 8'h2b;
	ram[820] = 8'hdf;	ram[821] = 8'hc2;	ram[822] = 8'h41;	ram[823] = 8'h03;
	ram[824] = 8'hdf;	ram[825] = 8'hcd;	ram[826] = 8'h8a;	ram[827] = 8'h05;
	ram[828] = 8'h21;	ram[829] = 8'h13;	ram[830] = 8'h01;	ram[831] = 8'h06;
	ram[832] = 8'h01;	ram[833] = 8'hcd;	ram[834] = 8'h82;	ram[835] = 8'h03;
	ram[836] = 8'hfe;	ram[837] = 8'h0d;	ram[838] = 8'hca;	ram[839] = 8'h85;
	ram[840] = 8'h05;	ram[841] = 8'hfe;	ram[842] = 8'h20;	ram[843] = 8'hda;
	ram[844] = 8'h41;	ram[845] = 8'h03;	ram[846] = 8'hfe;	ram[847] = 8'h7d;
	ram[848] = 8'hd2;	ram[849] = 8'h41;	ram[850] = 8'h03;	ram[851] = 8'hfe;
	ram[852] = 8'h40;	ram[853] = 8'hca;	ram[854] = 8'h38;	ram[855] = 8'h03;
	ram[856] = 8'hfe;	ram[857] = 8'h5f;	ram[858] = 8'hca;	ram[859] = 8'h32;
	ram[860] = 8'h03;	ram[861] = 8'h4f;	ram[862] = 8'h78;	ram[863] = 8'hfe;
	ram[864] = 8'h48;	ram[865] = 8'h3e;	ram[866] = 8'h07;	ram[867] = 8'hd2;
	ram[868] = 8'h6a;	ram[869] = 8'h03;	ram[870] = 8'h79;	ram[871] = 8'h71;
	ram[872] = 8'h23;	ram[873] = 8'h04;	ram[874] = 8'hdf;	ram[875] = 8'hc3;
	ram[876] = 8'h41;	ram[877] = 8'h03;	ram[878] = 8'hfe;	ram[879] = 8'h48;
	ram[880] = 8'hcc;	ram[881] = 8'h8a;	ram[882] = 8'h05;	ram[883] = 8'h3c;
	ram[884] = 8'h32;	ram[885] = 8'h27;	ram[886] = 8'h00;	ram[887] = 8'hdb;
	ram[888] = 8'h00;	ram[889] = 8'he6;	ram[890] = 8'h80;	ram[891] = 8'hc2;
	ram[892] = 8'h77;	ram[893] = 8'h03;	ram[894] = 8'hf1;	ram[895] = 8'hd3;
	ram[896] = 8'h01;	ram[897] = 8'hc9;	ram[898] = 8'hdb;	ram[899] = 8'h00;
	ram[900] = 8'he6;	ram[901] = 8'h01;	ram[902] = 8'hc2;	ram[903] = 8'h82;
	ram[904] = 8'h03;	ram[905] = 8'hdb;	ram[906] = 8'h01;	ram[907] = 8'he6;
	ram[908] = 8'h7f;	ram[909] = 8'hc9;	ram[910] = 8'hcd;	ram[911] = 8'h9d;
	ram[912] = 8'h04;	ram[913] = 8'hc0;	ram[914] = 8'hc1;	ram[915] = 8'hcd;
	ram[916] = 8'h7d;	ram[917] = 8'h02;	ram[918] = 8'hc5;	ram[919] = 8'he1;
	ram[920] = 8'hf7;	ram[921] = 8'hc1;	ram[922] = 8'h78;	ram[923] = 8'hb1;
	ram[924] = 8'hca;	ram[925] = 8'hf9;	ram[926] = 8'h01;	ram[927] = 8'hcd;
	ram[928] = 8'h73;	ram[929] = 8'h04;	ram[930] = 8'hc5;	ram[931] = 8'hcd;
	ram[932] = 8'h8a;	ram[933] = 8'h05;	ram[934] = 8'hf7;	ram[935] = 8'he3;
	ram[936] = 8'hcd;	ram[937] = 8'h37;	ram[938] = 8'h0b;	ram[939] = 8'h3e;
	ram[940] = 8'h20;	ram[941] = 8'he1;	ram[942] = 8'hdf;	ram[943] = 8'h7e;
	ram[944] = 8'hb7;	ram[945] = 8'h23;	ram[946] = 8'hca;	ram[947] = 8'h97;
	ram[948] = 8'h03;	ram[949] = 8'hf2;	ram[950] = 8'hae;	ram[951] = 8'h03;
	ram[952] = 8'hd6;	ram[953] = 8'h7f;	ram[954] = 8'h4f;	ram[955] = 8'he5;
	ram[956] = 8'h11;	ram[957] = 8'h57;	ram[958] = 8'h00;	ram[959] = 8'hd5;
	ram[960] = 8'h1a;	ram[961] = 8'h13;	ram[962] = 8'hb7;	ram[963] = 8'hf2;
	ram[964] = 8'hc0;	ram[965] = 8'h03;	ram[966] = 8'h0d;	ram[967] = 8'he1;
	ram[968] = 8'hc2;	ram[969] = 8'hbf;	ram[970] = 8'h03;	ram[971] = 8'h7e;
	ram[972] = 8'hb7;	ram[973] = 8'hfa;	ram[974] = 8'had;	ram[975] = 8'h03;
	ram[976] = 8'hdf;	ram[977] = 8'h23;	ram[978] = 8'hc3;	ram[979] = 8'hcb;
	ram[980] = 8'h03;	ram[981] = 8'hcd;	ram[982] = 8'h02;	ram[983] = 8'h05;
	ram[984] = 8'he3;	ram[985] = 8'hcd;	ram[986] = 8'h92;	ram[987] = 8'h01;
	ram[988] = 8'hd1;	ram[989] = 8'hc2;	ram[990] = 8'he2;	ram[991] = 8'h03;
	ram[992] = 8'h09;	ram[993] = 8'hf9;	ram[994] = 8'heb;	ram[995] = 8'h0e;
	ram[996] = 8'h08;	ram[997] = 8'hcd;	ram[998] = 8'hb6;	ram[999] = 8'h01;
	ram[1000] = 8'he5;	ram[1001] = 8'hcd;	ram[1002] = 8'hf5;	ram[1003] = 8'h04;
	ram[1004] = 8'he3;	ram[1005] = 8'he5;	ram[1006] = 8'h2a;	ram[1007] = 8'h61;
	ram[1008] = 8'h01;	ram[1009] = 8'he3;	ram[1010] = 8'hcf;	ram[1011] = 8'h95;
	ram[1012] = 8'hcd;	ram[1013] = 8'h8a;	ram[1014] = 8'h06;	ram[1015] = 8'he5;
	ram[1016] = 8'hcd;	ram[1017] = 8'h1d;	ram[1018] = 8'h0a;	ram[1019] = 8'he1;
	ram[1020] = 8'hc5;	ram[1021] = 8'hd5;	ram[1022] = 8'h01;	ram[1023] = 8'h00;
	ram[1024] = 8'h81;	ram[1025] = 8'h51;	ram[1026] = 8'h5a;	ram[1027] = 8'h7e;
	ram[1028] = 8'hfe;	ram[1029] = 8'h97;	ram[1030] = 8'h3e;	ram[1031] = 8'h01;
	ram[1032] = 8'hc2;	ram[1033] = 8'h14;	ram[1034] = 8'h04;	ram[1035] = 8'hcd;
	ram[1036] = 8'h8b;	ram[1037] = 8'h06;	ram[1038] = 8'he5;	ram[1039] = 8'hcd;
	ram[1040] = 8'h1d;	ram[1041] = 8'h0a;	ram[1042] = 8'hef;	ram[1043] = 8'he1;
	ram[1044] = 8'hc5;	ram[1045] = 8'hd5;	ram[1046] = 8'hf5;	ram[1047] = 8'h33;
	ram[1048] = 8'he5;	ram[1049] = 8'h2a;	ram[1050] = 8'h5d;	ram[1051] = 8'h01;
	ram[1052] = 8'he3;	ram[1053] = 8'h06;	ram[1054] = 8'h81;	ram[1055] = 8'hc5;
	ram[1056] = 8'h33;	ram[1057] = 8'hcd;	ram[1058] = 8'h73;	ram[1059] = 8'h04;
	ram[1060] = 8'h7e;	ram[1061] = 8'hfe;	ram[1062] = 8'h3a;	ram[1063] = 8'hca;
	ram[1064] = 8'h3e;	ram[1065] = 8'h04;	ram[1066] = 8'hb7;	ram[1067] = 8'hc2;
	ram[1068] = 8'hd0;	ram[1069] = 8'h01;	ram[1070] = 8'h23;	ram[1071] = 8'h7e;
	ram[1072] = 8'h23;	ram[1073] = 8'hb6;	ram[1074] = 8'h23;	ram[1075] = 8'hca;
	ram[1076] = 8'hf9;	ram[1077] = 8'h01;	ram[1078] = 8'h5e;	ram[1079] = 8'h23;
	ram[1080] = 8'h56;	ram[1081] = 8'heb;	ram[1082] = 8'h22;	ram[1083] = 8'h61;
	ram[1084] = 8'h01;	ram[1085] = 8'heb;	ram[1086] = 8'hd7;	ram[1087] = 8'h11;
	ram[1088] = 8'h21;	ram[1089] = 8'h04;	ram[1090] = 8'hd5;	ram[1091] = 8'hc8;
	ram[1092] = 8'hd6;	ram[1093] = 8'h80;	ram[1094] = 8'hda;	ram[1095] = 8'h02;
	ram[1096] = 8'h05;	ram[1097] = 8'hfe;	ram[1098] = 8'h14;	ram[1099] = 8'hd2;
	ram[1100] = 8'hd0;	ram[1101] = 8'h01;	ram[1102] = 8'h07;	ram[1103] = 8'h4f;
	ram[1104] = 8'h06;	ram[1105] = 8'h00;	ram[1106] = 8'heb;	ram[1107] = 8'h21;
	ram[1108] = 8'hd2;	ram[1109] = 8'h00;	ram[1110] = 8'h09;	ram[1111] = 8'h4e;
	ram[1112] = 8'h23;	ram[1113] = 8'h46;	ram[1114] = 8'hc5;	ram[1115] = 8'heb;
	ram[1116] = 8'hd7;	ram[1117] = 8'hc9;	ram[1118] = 8'hfe;	ram[1119] = 8'h20;
	ram[1120] = 8'hca;	ram[1121] = 8'h10;	ram[1122] = 8'h00;	ram[1123] = 8'hfe;
	ram[1124] = 8'h30;	ram[1125] = 8'h3f;	ram[1126] = 8'h3c;	ram[1127] = 8'h3d;
	ram[1128] = 8'hc9;	ram[1129] = 8'heb;	ram[1130] = 8'h2a;	ram[1131] = 8'h65;
	ram[1132] = 8'h01;	ram[1133] = 8'h2b;	ram[1134] = 8'h22;	ram[1135] = 8'h6d;
	ram[1136] = 8'h01;	ram[1137] = 8'heb;	ram[1138] = 8'hc9;	ram[1139] = 8'hdb;
	ram[1140] = 8'h00;	ram[1141] = 8'he6;	ram[1142] = 8'h01;	ram[1143] = 8'hc0;
	ram[1144] = 8'hcd;	ram[1145] = 8'h82;	ram[1146] = 8'h03;	ram[1147] = 8'hfe;
	ram[1148] = 8'h03;	ram[1149] = 8'hc3;	ram[1150] = 8'hf7;	ram[1151] = 8'h01;
	ram[1152] = 8'h7e;	ram[1153] = 8'hfe;	ram[1154] = 8'h41;	ram[1155] = 8'hd8;
	ram[1156] = 8'hfe;	ram[1157] = 8'h5b;	ram[1158] = 8'h3f;	ram[1159] = 8'hc9;
	ram[1160] = 8'hd7;	ram[1161] = 8'hcd;	ram[1162] = 8'h8a;	ram[1163] = 8'h06;
	ram[1164] = 8'hef;	ram[1165] = 8'hfa;	ram[1166] = 8'h98;	ram[1167] = 8'h04;
	ram[1168] = 8'h3a;	ram[1169] = 8'h72;	ram[1170] = 8'h01;	ram[1171] = 8'hfe;
	ram[1172] = 8'h90;	ram[1173] = 8'hda;	ram[1174] = 8'h77;	ram[1175] = 8'h0a;
	ram[1176] = 8'h1e;	ram[1177] = 8'h08;	ram[1178] = 8'hc3;	ram[1179] = 8'hd5;
	ram[1180] = 8'h01;	ram[1181] = 8'h2b;	ram[1182] = 8'h11;	ram[1183] = 8'h00;
	ram[1184] = 8'h00;	ram[1185] = 8'hd7;	ram[1186] = 8'hd0;	ram[1187] = 8'he5;
	ram[1188] = 8'hf5;	ram[1189] = 8'h21;	ram[1190] = 8'h98;	ram[1191] = 8'h19;
	ram[1192] = 8'he7;	ram[1193] = 8'hda;	ram[1194] = 8'hd0;	ram[1195] = 8'h01;
	ram[1196] = 8'h62;	ram[1197] = 8'h6b;	ram[1198] = 8'h19;	ram[1199] = 8'h29;
	ram[1200] = 8'h19;	ram[1201] = 8'h29;	ram[1202] = 8'hf1;	ram[1203] = 8'hd6;
	ram[1204] = 8'h30;	ram[1205] = 8'h5f;	ram[1206] = 8'h16;	ram[1207] = 8'h00;
	ram[1208] = 8'h19;	ram[1209] = 8'heb;	ram[1210] = 8'he1;	ram[1211] = 8'hc3;
	ram[1212] = 8'ha1;	ram[1213] = 8'h04;	ram[1214] = 8'h0e;	ram[1215] = 8'h03;
	ram[1216] = 8'hcd;	ram[1217] = 8'hb6;	ram[1218] = 8'h01;	ram[1219] = 8'hc1;
	ram[1220] = 8'he5;	ram[1221] = 8'he5;	ram[1222] = 8'h2a;	ram[1223] = 8'h61;
	ram[1224] = 8'h01;	ram[1225] = 8'he3;	ram[1226] = 8'h16;	ram[1227] = 8'h8c;
	ram[1228] = 8'hd5;	ram[1229] = 8'h33;	ram[1230] = 8'hc5;	ram[1231] = 8'hcd;
	ram[1232] = 8'h9d;	ram[1233] = 8'h04;	ram[1234] = 8'hc0;	ram[1235] = 8'hcd;
	ram[1236] = 8'h7d;	ram[1237] = 8'h02;	ram[1238] = 8'h60;	ram[1239] = 8'h69;
	ram[1240] = 8'h2b;	ram[1241] = 8'hd8;	ram[1242] = 8'h1e;	ram[1243] = 8'h0e;
	ram[1244] = 8'hc3;	ram[1245] = 8'hd5;	ram[1246] = 8'h01;	ram[1247] = 8'hc0;
	ram[1248] = 8'h16;	ram[1249] = 8'hff;	ram[1250] = 8'hcd;	ram[1251] = 8'h92;
	ram[1252] = 8'h01;	ram[1253] = 8'hf9;	ram[1254] = 8'hfe;	ram[1255] = 8'h8c;
	ram[1256] = 8'h1e;	ram[1257] = 8'h04;	ram[1258] = 8'hc2;	ram[1259] = 8'hd5;
	ram[1260] = 8'h01;	ram[1261] = 8'he1;	ram[1262] = 8'h22;	ram[1263] = 8'h61;
	ram[1264] = 8'h01;	ram[1265] = 8'h21;	ram[1266] = 8'h21;	ram[1267] = 8'h04;
	ram[1268] = 8'he3;	ram[1269] = 8'h01;	ram[1270] = 8'h3a;	ram[1271] = 8'h10;
	ram[1272] = 8'h00;	ram[1273] = 8'h7e;	ram[1274] = 8'hb7;	ram[1275] = 8'hc8;
	ram[1276] = 8'hb9;	ram[1277] = 8'hc8;	ram[1278] = 8'h23;	ram[1279] = 8'hc3;
	ram[1280] = 8'hf9;	ram[1281] = 8'h04;	ram[1282] = 8'hcd;	ram[1283] = 8'h1b;
	ram[1284] = 8'h07;	ram[1285] = 8'hcf;	ram[1286] = 8'h9d;	ram[1287] = 8'hd5;
	ram[1288] = 8'hcd;	ram[1289] = 8'h8a;	ram[1290] = 8'h06;	ram[1291] = 8'he3;
	ram[1292] = 8'h22;	ram[1293] = 8'h5d;	ram[1294] = 8'h01;	ram[1295] = 8'he5;
	ram[1296] = 8'hcd;	ram[1297] = 8'h29;	ram[1298] = 8'h0a;	ram[1299] = 8'hd1;
	ram[1300] = 8'he1;	ram[1301] = 8'hc9;	ram[1302] = 8'hcd;	ram[1303] = 8'h8a;
	ram[1304] = 8'h06;	ram[1305] = 8'h7e;	ram[1306] = 8'hcd;	ram[1307] = 8'h02;
	ram[1308] = 8'h0a;	ram[1309] = 8'h16;	ram[1310] = 8'h00;	ram[1311] = 8'hd6;
	ram[1312] = 8'h9c;	ram[1313] = 8'hda;	ram[1314] = 8'h32;	ram[1315] = 8'h05;
	ram[1316] = 8'hfe;	ram[1317] = 8'h03;	ram[1318] = 8'hd2;	ram[1319] = 8'h32;
	ram[1320] = 8'h05;	ram[1321] = 8'hfe;	ram[1322] = 8'h01;	ram[1323] = 8'h17;
	ram[1324] = 8'hb2;	ram[1325] = 8'h57;	ram[1326] = 8'hd7;	ram[1327] = 8'hc3;
	ram[1328] = 8'h1f;	ram[1329] = 8'h05;	ram[1330] = 8'h7a;	ram[1331] = 8'hb7;
	ram[1332] = 8'hca;	ram[1333] = 8'hd0;	ram[1334] = 8'h01;	ram[1335] = 8'hf5;
	ram[1336] = 8'hcd;	ram[1337] = 8'h8a;	ram[1338] = 8'h06;	ram[1339] = 8'hcf;
	ram[1340] = 8'h96;	ram[1341] = 8'h2b;	ram[1342] = 8'hf1;	ram[1343] = 8'hc1;
	ram[1344] = 8'hd1;	ram[1345] = 8'he5;	ram[1346] = 8'hf5;	ram[1347] = 8'hcd;
	ram[1348] = 8'h4c;	ram[1349] = 8'h0a;	ram[1350] = 8'h3c;	ram[1351] = 8'h17;
	ram[1352] = 8'hc1;	ram[1353] = 8'ha0;	ram[1354] = 8'he1;	ram[1355] = 8'hca;
	ram[1356] = 8'hf7;	ram[1357] = 8'h04;	ram[1358] = 8'hd7;	ram[1359] = 8'hda;
	ram[1360] = 8'hcf;	ram[1361] = 8'h04;	ram[1362] = 8'hc3;	ram[1363] = 8'h43;
	ram[1364] = 8'h04;	ram[1365] = 8'h2b;	ram[1366] = 8'hd7;	ram[1367] = 8'hca;
	ram[1368] = 8'h8a;	ram[1369] = 8'h05;	ram[1370] = 8'hc8;	ram[1371] = 8'hfe;
	ram[1372] = 8'h22;	ram[1373] = 8'hcc;	ram[1374] = 8'ha2;	ram[1375] = 8'h05;
	ram[1376] = 8'hca;	ram[1377] = 8'h55;	ram[1378] = 8'h05;	ram[1379] = 8'hfe;
	ram[1380] = 8'h94;	ram[1381] = 8'hca;	ram[1382] = 8'hc7;	ram[1383] = 8'h05;
	ram[1384] = 8'he5;	ram[1385] = 8'hfe;	ram[1386] = 8'h2c;	ram[1387] = 8'hca;
	ram[1388] = 8'hb3;	ram[1389] = 8'h05;	ram[1390] = 8'hfe;	ram[1391] = 8'h3b;
	ram[1392] = 8'hca;	ram[1393] = 8'hdf;	ram[1394] = 8'h05;	ram[1395] = 8'hc1;
	ram[1396] = 8'hcd;	ram[1397] = 8'h8a;	ram[1398] = 8'h06;	ram[1399] = 8'he5;
	ram[1400] = 8'hcd;	ram[1401] = 8'h42;	ram[1402] = 8'h0b;	ram[1403] = 8'hcd;
	ram[1404] = 8'ha3;	ram[1405] = 8'h05;	ram[1406] = 8'h3e;	ram[1407] = 8'h20;
	ram[1408] = 8'hdf;	ram[1409] = 8'he1;	ram[1410] = 8'hc3;	ram[1411] = 8'h55;
	ram[1412] = 8'h05;	ram[1413] = 8'h36;	ram[1414] = 8'h00;	ram[1415] = 8'h21;
	ram[1416] = 8'h12;	ram[1417] = 8'h01;	ram[1418] = 8'h3e;	ram[1419] = 8'h0d;
	ram[1420] = 8'h32;	ram[1421] = 8'h27;	ram[1422] = 8'h00;	ram[1423] = 8'hdf;
	ram[1424] = 8'h3e;	ram[1425] = 8'h0a;	ram[1426] = 8'hdf;	ram[1427] = 8'h3a;
	ram[1428] = 8'h26;	ram[1429] = 8'h00;	ram[1430] = 8'h3d;	ram[1431] = 8'h32;
	ram[1432] = 8'h27;	ram[1433] = 8'h00;	ram[1434] = 8'hc8;	ram[1435] = 8'hf5;
	ram[1436] = 8'haf;	ram[1437] = 8'hdf;	ram[1438] = 8'hf1;	ram[1439] = 8'hc3;
	ram[1440] = 8'h96;	ram[1441] = 8'h05;	ram[1442] = 8'h23;	ram[1443] = 8'h7e;
	ram[1444] = 8'hb7;	ram[1445] = 8'hc8;	ram[1446] = 8'h23;	ram[1447] = 8'hfe;
	ram[1448] = 8'h22;	ram[1449] = 8'hc8;	ram[1450] = 8'hdf;	ram[1451] = 8'hfe;
	ram[1452] = 8'h0d;	ram[1453] = 8'hcc;	ram[1454] = 8'h8a;	ram[1455] = 8'h05;
	ram[1456] = 8'hc3;	ram[1457] = 8'ha3;	ram[1458] = 8'h05;	ram[1459] = 8'h3a;
	ram[1460] = 8'h27;	ram[1461] = 8'h00;	ram[1462] = 8'hfe;	ram[1463] = 8'h38;
	ram[1464] = 8'hd4;	ram[1465] = 8'h8a;	ram[1466] = 8'h05;	ram[1467] = 8'hd2;
	ram[1468] = 8'hdf;	ram[1469] = 8'h05;	ram[1470] = 8'hd6;	ram[1471] = 8'h0e;
	ram[1472] = 8'hd2;	ram[1473] = 8'hbe;	ram[1474] = 8'h05;	ram[1475] = 8'h2f;
	ram[1476] = 8'hc3;	ram[1477] = 8'hd6;	ram[1478] = 8'h05;	ram[1479] = 8'hcd;
	ram[1480] = 8'h88;	ram[1481] = 8'h04;	ram[1482] = 8'hcf;	ram[1483] = 8'h29;
	ram[1484] = 8'h2b;	ram[1485] = 8'he5;	ram[1486] = 8'h3a;	ram[1487] = 8'h27;
	ram[1488] = 8'h00;	ram[1489] = 8'h2f;	ram[1490] = 8'h83;	ram[1491] = 8'hd2;
	ram[1492] = 8'hdf;	ram[1493] = 8'h05;	ram[1494] = 8'h3c;	ram[1495] = 8'h47;
	ram[1496] = 8'h3e;	ram[1497] = 8'h20;	ram[1498] = 8'hdf;	ram[1499] = 8'h05;
	ram[1500] = 8'hc2;	ram[1501] = 8'hda;	ram[1502] = 8'h05;	ram[1503] = 8'he1;
	ram[1504] = 8'hd7;	ram[1505] = 8'hc3;	ram[1506] = 8'h5a;	ram[1507] = 8'h05;
	ram[1508] = 8'he5;	ram[1509] = 8'h2a;	ram[1510] = 8'h61;	ram[1511] = 8'h01;
	ram[1512] = 8'h1e;	ram[1513] = 8'h16;	ram[1514] = 8'h23;	ram[1515] = 8'h7d;
	ram[1516] = 8'hb4;	ram[1517] = 8'hca;	ram[1518] = 8'hd5;	ram[1519] = 8'h01;
	ram[1520] = 8'hcd;	ram[1521] = 8'hc2;	ram[1522] = 8'h02;	ram[1523] = 8'hc3;
	ram[1524] = 8'hfb;	ram[1525] = 8'h05;	ram[1526] = 8'he5;	ram[1527] = 8'h2a;
	ram[1528] = 8'h6d;	ram[1529] = 8'h01;	ram[1530] = 8'hf6;	ram[1531] = 8'haf;
	ram[1532] = 8'h32;	ram[1533] = 8'h5c;	ram[1534] = 8'h01;	ram[1535] = 8'he3;
	ram[1536] = 8'h01;	ram[1537] = 8'hcf;	ram[1538] = 8'h2c;	ram[1539] = 8'hcd;
	ram[1540] = 8'h1b;	ram[1541] = 8'h07;	ram[1542] = 8'he3;	ram[1543] = 8'hd5;
	ram[1544] = 8'h7e;	ram[1545] = 8'hfe;	ram[1546] = 8'h2c;	ram[1547] = 8'hca;
	ram[1548] = 8'h20;	ram[1549] = 8'h06;	ram[1550] = 8'hb7;	ram[1551] = 8'hc2;
	ram[1552] = 8'hd0;	ram[1553] = 8'h01;	ram[1554] = 8'h3a;	ram[1555] = 8'h5c;
	ram[1556] = 8'h01;	ram[1557] = 8'hb7;	ram[1558] = 8'h23;	ram[1559] = 8'hc2;
	ram[1560] = 8'h36;	ram[1561] = 8'h06;	ram[1562] = 8'h3e;	ram[1563] = 8'h3f;
	ram[1564] = 8'hdf;	ram[1565] = 8'hcd;	ram[1566] = 8'hc2;	ram[1567] = 8'h02;
	ram[1568] = 8'hd1;	ram[1569] = 8'h23;	ram[1570] = 8'hcd;	ram[1571] = 8'h07;
	ram[1572] = 8'h05;	ram[1573] = 8'he3;	ram[1574] = 8'h2b;	ram[1575] = 8'hd7;
	ram[1576] = 8'hc2;	ram[1577] = 8'h01;	ram[1578] = 8'h06;	ram[1579] = 8'hd1;
	ram[1580] = 8'h3a;	ram[1581] = 8'h5c;	ram[1582] = 8'h01;	ram[1583] = 8'hb7;
	ram[1584] = 8'hc8;	ram[1585] = 8'heb;	ram[1586] = 8'hc2;	ram[1587] = 8'h6e;
	ram[1588] = 8'h04;	ram[1589] = 8'he1;	ram[1590] = 8'hf7;	ram[1591] = 8'h79;
	ram[1592] = 8'hb0;	ram[1593] = 8'h1e;	ram[1594] = 8'h06;	ram[1595] = 8'hca;
	ram[1596] = 8'hd5;	ram[1597] = 8'h01;	ram[1598] = 8'h23;	ram[1599] = 8'hd7;
	ram[1600] = 8'hfe;	ram[1601] = 8'h83;	ram[1602] = 8'hc2;	ram[1603] = 8'h35;
	ram[1604] = 8'h06;	ram[1605] = 8'hc1;	ram[1606] = 8'hc3;	ram[1607] = 8'h20;
	ram[1608] = 8'h06;	ram[1609] = 8'hcd;	ram[1610] = 8'h1b;	ram[1611] = 8'h07;
	ram[1612] = 8'h22;	ram[1613] = 8'h5d;	ram[1614] = 8'h01;	ram[1615] = 8'hcd;
	ram[1616] = 8'h92;	ram[1617] = 8'h01;	ram[1618] = 8'hf9;	ram[1619] = 8'hd5;
	ram[1620] = 8'h7e;	ram[1621] = 8'h23;	ram[1622] = 8'hf5;	ram[1623] = 8'hd5;
	ram[1624] = 8'h1e;	ram[1625] = 8'h00;	ram[1626] = 8'hc2;	ram[1627] = 8'hd5;
	ram[1628] = 8'h01;	ram[1629] = 8'hcd;	ram[1630] = 8'h0f;	ram[1631] = 8'h0a;
	ram[1632] = 8'he3;	ram[1633] = 8'he5;	ram[1634] = 8'hcd;	ram[1635] = 8'h04;
	ram[1636] = 8'h08;	ram[1637] = 8'he1;	ram[1638] = 8'hcd;	ram[1639] = 8'h29;
	ram[1640] = 8'h0a;	ram[1641] = 8'he1;	ram[1642] = 8'hcd;	ram[1643] = 8'h20;
	ram[1644] = 8'h0a;	ram[1645] = 8'he5;	ram[1646] = 8'hcd;	ram[1647] = 8'h4c;
	ram[1648] = 8'h0a;	ram[1649] = 8'he1;	ram[1650] = 8'hc1;	ram[1651] = 8'h90;
	ram[1652] = 8'hcd;	ram[1653] = 8'h20;	ram[1654] = 8'h0a;	ram[1655] = 8'hca;
	ram[1656] = 8'h83;	ram[1657] = 8'h06;	ram[1658] = 8'heb;	ram[1659] = 8'h22;
	ram[1660] = 8'h61;	ram[1661] = 8'h01;	ram[1662] = 8'h69;	ram[1663] = 8'h60;
	ram[1664] = 8'hc3;	ram[1665] = 8'h1d;	ram[1666] = 8'h04;	ram[1667] = 8'hf9;
	ram[1668] = 8'h2a;	ram[1669] = 8'h5d;	ram[1670] = 8'h01;	ram[1671] = 8'hc3;
	ram[1672] = 8'h21;	ram[1673] = 8'h04;	ram[1674] = 8'h2b;	ram[1675] = 8'h16;
	ram[1676] = 8'h00;	ram[1677] = 8'hd5;	ram[1678] = 8'h0e;	ram[1679] = 8'h01;
	ram[1680] = 8'hcd;	ram[1681] = 8'hb6;	ram[1682] = 8'h01;	ram[1683] = 8'hcd;
	ram[1684] = 8'hc4;	ram[1685] = 8'h06;	ram[1686] = 8'h22;	ram[1687] = 8'h5f;
	ram[1688] = 8'h01;	ram[1689] = 8'h2a;	ram[1690] = 8'h5f;	ram[1691] = 8'h01;
	ram[1692] = 8'hc1;	ram[1693] = 8'h7e;	ram[1694] = 8'h16;	ram[1695] = 8'h00;
	ram[1696] = 8'hd6;	ram[1697] = 8'h98;	ram[1698] = 8'hd8;	ram[1699] = 8'hfe;
	ram[1700] = 8'h04;	ram[1701] = 8'hd0;	ram[1702] = 8'h5f;	ram[1703] = 8'h07;
	ram[1704] = 8'h83;	ram[1705] = 8'h5f;	ram[1706] = 8'h21;	ram[1707] = 8'h4b;
	ram[1708] = 8'h00;	ram[1709] = 8'h19;	ram[1710] = 8'h78;	ram[1711] = 8'h56;
	ram[1712] = 8'hba;	ram[1713] = 8'hd0;	ram[1714] = 8'h23;	ram[1715] = 8'hc5;
	ram[1716] = 8'h01;	ram[1717] = 8'h99;	ram[1718] = 8'h06;	ram[1719] = 8'hc5;
	ram[1720] = 8'h4a;	ram[1721] = 8'hcd;	ram[1722] = 8'h02;	ram[1723] = 8'h0a;
	ram[1724] = 8'h51;	ram[1725] = 8'hf7;	ram[1726] = 8'h2a;	ram[1727] = 8'h5f;
	ram[1728] = 8'h01;	ram[1729] = 8'hc3;	ram[1730] = 8'h8d;	ram[1731] = 8'h06;
	ram[1732] = 8'hd7;	ram[1733] = 8'hda;	ram[1734] = 8'hb3;	ram[1735] = 8'h0a;
	ram[1736] = 8'hcd;	ram[1737] = 8'h80;	ram[1738] = 8'h04;	ram[1739] = 8'hd2;
	ram[1740] = 8'hf3;	ram[1741] = 8'h06;	ram[1742] = 8'hfe;	ram[1743] = 8'h98;
	ram[1744] = 8'hca;	ram[1745] = 8'hc4;	ram[1746] = 8'h06;	ram[1747] = 8'hfe;
	ram[1748] = 8'h2e;	ram[1749] = 8'hca;	ram[1750] = 8'hb3;	ram[1751] = 8'h0a;
	ram[1752] = 8'hfe;	ram[1753] = 8'h99;	ram[1754] = 8'hca;	ram[1755] = 8'hea;
	ram[1756] = 8'h06;	ram[1757] = 8'hd6;	ram[1758] = 8'h9f;	ram[1759] = 8'hd2;
	ram[1760] = 8'hfd;	ram[1761] = 8'h06;	ram[1762] = 8'hcf;	ram[1763] = 8'h28;
	ram[1764] = 8'hcd;	ram[1765] = 8'h8a;	ram[1766] = 8'h06;	ram[1767] = 8'hcf;
	ram[1768] = 8'h29;	ram[1769] = 8'hc9;	ram[1770] = 8'hcd;	ram[1771] = 8'hc4;
	ram[1772] = 8'h06;	ram[1773] = 8'he5;	ram[1774] = 8'hcd;	ram[1775] = 8'hfa;
	ram[1776] = 8'h09;	ram[1777] = 8'he1;	ram[1778] = 8'hc9;	ram[1779] = 8'hcd;
	ram[1780] = 8'h1b;	ram[1781] = 8'h07;	ram[1782] = 8'he5;	ram[1783] = 8'heb;
	ram[1784] = 8'hcd;	ram[1785] = 8'h0f;	ram[1786] = 8'h0a;	ram[1787] = 8'he1;
	ram[1788] = 8'hc9;	ram[1789] = 8'h06;	ram[1790] = 8'h00;	ram[1791] = 8'h07;
	ram[1792] = 8'h4f;	ram[1793] = 8'hc5;	ram[1794] = 8'hd7;	ram[1795] = 8'hcd;
	ram[1796] = 8'he2;	ram[1797] = 8'h06;	ram[1798] = 8'he3;	ram[1799] = 8'h11;
	ram[1800] = 8'hf1;	ram[1801] = 8'h06;	ram[1802] = 8'hd5;	ram[1803] = 8'h01;
	ram[1804] = 8'h3d;	ram[1805] = 8'h00;	ram[1806] = 8'h09;	ram[1807] = 8'hf7;
	ram[1808] = 8'hc9;	ram[1809] = 8'h2b;	ram[1810] = 8'hd7;	ram[1811] = 8'hc8;
	ram[1812] = 8'hcf;	ram[1813] = 8'h2c;	ram[1814] = 8'h01;	ram[1815] = 8'h11;
	ram[1816] = 8'h07;	ram[1817] = 8'hc5;	ram[1818] = 8'hf6;	ram[1819] = 8'haf;
	ram[1820] = 8'h32;	ram[1821] = 8'h5b;	ram[1822] = 8'h01;	ram[1823] = 8'h46;
	ram[1824] = 8'hcd;	ram[1825] = 8'h80;	ram[1826] = 8'h04;	ram[1827] = 8'hda;
	ram[1828] = 8'hd0;	ram[1829] = 8'h01;	ram[1830] = 8'haf;	ram[1831] = 8'h4f;
	ram[1832] = 8'hd7;	ram[1833] = 8'hd2;	ram[1834] = 8'h2e;	ram[1835] = 8'h07;
	ram[1836] = 8'h4f;	ram[1837] = 8'hd7;	ram[1838] = 8'hd6;	ram[1839] = 8'h28;
	ram[1840] = 8'hca;	ram[1841] = 8'h8a;	ram[1842] = 8'h07;	ram[1843] = 8'he5;
	ram[1844] = 8'h2a;	ram[1845] = 8'h69;	ram[1846] = 8'h01;	ram[1847] = 8'heb;
	ram[1848] = 8'h2a;	ram[1849] = 8'h67;	ram[1850] = 8'h01;	ram[1851] = 8'he7;
	ram[1852] = 8'hca;	ram[1853] = 8'h52;	ram[1854] = 8'h07;	ram[1855] = 8'h79;
	ram[1856] = 8'h96;	ram[1857] = 8'h23;	ram[1858] = 8'hc2;	ram[1859] = 8'h47;
	ram[1860] = 8'h07;	ram[1861] = 8'h78;	ram[1862] = 8'h96;	ram[1863] = 8'h23;
	ram[1864] = 8'hca;	ram[1865] = 8'h82;	ram[1866] = 8'h07;	ram[1867] = 8'h23;
	ram[1868] = 8'h23;	ram[1869] = 8'h23;	ram[1870] = 8'h23;	ram[1871] = 8'hc3;
	ram[1872] = 8'h3b;	ram[1873] = 8'h07;	ram[1874] = 8'he1;	ram[1875] = 8'he3;
	ram[1876] = 8'hd5;	ram[1877] = 8'h11;	ram[1878] = 8'hf6;	ram[1879] = 8'h06;
	ram[1880] = 8'he7;	ram[1881] = 8'hd1;	ram[1882] = 8'hca;	ram[1883] = 8'h85;
	ram[1884] = 8'h07;	ram[1885] = 8'he3;	ram[1886] = 8'he5;	ram[1887] = 8'hc5;
	ram[1888] = 8'h01;	ram[1889] = 8'h06;	ram[1890] = 8'h00;	ram[1891] = 8'h2a;
	ram[1892] = 8'h6b;	ram[1893] = 8'h01;	ram[1894] = 8'he5;	ram[1895] = 8'h09;
	ram[1896] = 8'hc1;	ram[1897] = 8'he5;	ram[1898] = 8'hcd;	ram[1899] = 8'ha7;
	ram[1900] = 8'h01;	ram[1901] = 8'he1;	ram[1902] = 8'h22;	ram[1903] = 8'h6b;
	ram[1904] = 8'h01;	ram[1905] = 8'h60;	ram[1906] = 8'h69;	ram[1907] = 8'h22;
	ram[1908] = 8'h69;	ram[1909] = 8'h01;	ram[1910] = 8'h2b;	ram[1911] = 8'h36;
	ram[1912] = 8'h00;	ram[1913] = 8'he7;	ram[1914] = 8'hc2;	ram[1915] = 8'h76;
	ram[1916] = 8'h07;	ram[1917] = 8'hd1;	ram[1918] = 8'h73;	ram[1919] = 8'h23;
	ram[1920] = 8'h72;	ram[1921] = 8'h23;	ram[1922] = 8'heb;	ram[1923] = 8'he1;
	ram[1924] = 8'hc9;	ram[1925] = 8'h32;	ram[1926] = 8'h72;	ram[1927] = 8'h01;
	ram[1928] = 8'he1;	ram[1929] = 8'hc9;	ram[1930] = 8'hc5;	ram[1931] = 8'h3a;
	ram[1932] = 8'h5b;	ram[1933] = 8'h01;	ram[1934] = 8'hf5;	ram[1935] = 8'hcd;
	ram[1936] = 8'h88;	ram[1937] = 8'h04;	ram[1938] = 8'hcf;	ram[1939] = 8'h29;
	ram[1940] = 8'hf1;	ram[1941] = 8'h32;	ram[1942] = 8'h5b;	ram[1943] = 8'h01;
	ram[1944] = 8'he3;	ram[1945] = 8'heb;	ram[1946] = 8'h29;	ram[1947] = 8'h29;
	ram[1948] = 8'he5;	ram[1949] = 8'h2a;	ram[1950] = 8'h69;	ram[1951] = 8'h01;
	ram[1952] = 8'h01;	ram[1953] = 8'hc1;	ram[1954] = 8'h09;	ram[1955] = 8'heb;
	ram[1956] = 8'he5;	ram[1957] = 8'h2a;	ram[1958] = 8'h6b;	ram[1959] = 8'h01;
	ram[1960] = 8'he7;	ram[1961] = 8'heb;	ram[1962] = 8'hd1;	ram[1963] = 8'hca;
	ram[1964] = 8'hcd;	ram[1965] = 8'h07;	ram[1966] = 8'hf7;	ram[1967] = 8'he3;
	ram[1968] = 8'he7;	ram[1969] = 8'he1;	ram[1970] = 8'hf7;	ram[1971] = 8'hc2;
	ram[1972] = 8'ha1;	ram[1973] = 8'h07;	ram[1974] = 8'h3a;	ram[1975] = 8'h5b;
	ram[1976] = 8'h01;	ram[1977] = 8'hb7;	ram[1978] = 8'h1e;	ram[1979] = 8'h12;
	ram[1980] = 8'hc2;	ram[1981] = 8'hd5;	ram[1982] = 8'h01;	ram[1983] = 8'hd1;
	ram[1984] = 8'h1b;	ram[1985] = 8'he3;	ram[1986] = 8'he7;	ram[1987] = 8'h1e;
	ram[1988] = 8'h10;	ram[1989] = 8'hd2;	ram[1990] = 8'hd5;	ram[1991] = 8'h01;
	ram[1992] = 8'hd1;	ram[1993] = 8'h19;	ram[1994] = 8'hd1;	ram[1995] = 8'heb;
	ram[1996] = 8'hc9;	ram[1997] = 8'h73;	ram[1998] = 8'h23;	ram[1999] = 8'h72;
	ram[2000] = 8'h23;	ram[2001] = 8'h11;	ram[2002] = 8'h2c;	ram[2003] = 8'h00;
	ram[2004] = 8'h3a;	ram[2005] = 8'h5b;	ram[2006] = 8'h01;	ram[2007] = 8'hb7;
	ram[2008] = 8'hca;	ram[2009] = 8'he1;	ram[2010] = 8'h07;	ram[2011] = 8'hd1;
	ram[2012] = 8'hd5;	ram[2013] = 8'h13;	ram[2014] = 8'h13;	ram[2015] = 8'h13;
	ram[2016] = 8'h13;	ram[2017] = 8'hd5;	ram[2018] = 8'h73;	ram[2019] = 8'h23;
	ram[2020] = 8'h72;	ram[2021] = 8'h23;	ram[2022] = 8'he5;	ram[2023] = 8'h19;
	ram[2024] = 8'hcd;	ram[2025] = 8'hc3;	ram[2026] = 8'h01;	ram[2027] = 8'h22;
	ram[2028] = 8'h6b;	ram[2029] = 8'h01;	ram[2030] = 8'hd1;	ram[2031] = 8'h2b;
	ram[2032] = 8'h36;	ram[2033] = 8'h00;	ram[2034] = 8'he7;	ram[2035] = 8'hc2;
	ram[2036] = 8'hef;	ram[2037] = 8'h07;	ram[2038] = 8'hc3;	ram[2039] = 8'hbf;
	ram[2040] = 8'h07;	ram[2041] = 8'h50;	ram[2042] = 8'h1e;	ram[2043] = 8'h00;
	ram[2044] = 8'h06;	ram[2045] = 8'h90;	ram[2046] = 8'hc3;	ram[2047] = 8'hea;
	ram[2048] = 8'h09;	ram[2049] = 8'h21;	ram[2050] = 8'h0b;	ram[2051] = 8'h0c;
	ram[2052] = 8'hcd;	ram[2053] = 8'h20;	ram[2054] = 8'h0a;	ram[2055] = 8'hc3;
	ram[2056] = 8'h12;	ram[2057] = 8'h08;	ram[2058] = 8'hc1;	ram[2059] = 8'hd1;
	ram[2060] = 8'hcd;	ram[2061] = 8'hfa;	ram[2062] = 8'h09;	ram[2063] = 8'h21;
	ram[2064] = 8'hc1;	ram[2065] = 8'hd1;	ram[2066] = 8'h78;	ram[2067] = 8'hb7;
	ram[2068] = 8'hc8;	ram[2069] = 8'h3a;	ram[2070] = 8'h72;	ram[2071] = 8'h01;
	ram[2072] = 8'hb7;	ram[2073] = 8'hca;	ram[2074] = 8'h12;	ram[2075] = 8'h0a;
	ram[2076] = 8'h90;	ram[2077] = 8'hd2;	ram[2078] = 8'h2c;	ram[2079] = 8'h08;
	ram[2080] = 8'h2f;	ram[2081] = 8'h3c;	ram[2082] = 8'heb;	ram[2083] = 8'hcd;
	ram[2084] = 8'h02;	ram[2085] = 8'h0a;	ram[2086] = 8'heb;	ram[2087] = 8'hcd;
	ram[2088] = 8'h12;	ram[2089] = 8'h0a;	ram[2090] = 8'hc1;	ram[2091] = 8'hd1;
	ram[2092] = 8'hf5;	ram[2093] = 8'hcd;	ram[2094] = 8'h37;	ram[2095] = 8'h0a;
	ram[2096] = 8'h67;	ram[2097] = 8'hf1;	ram[2098] = 8'hcd;	ram[2099] = 8'hc9;
	ram[2100] = 8'h08;	ram[2101] = 8'hb4;	ram[2102] = 8'h21;	ram[2103] = 8'h6f;
	ram[2104] = 8'h01;	ram[2105] = 8'hf2;	ram[2106] = 8'h4d;	ram[2107] = 8'h08;
	ram[2108] = 8'hcd;	ram[2109] = 8'ha9;	ram[2110] = 8'h08;	ram[2111] = 8'hd2;
	ram[2112] = 8'h7e;	ram[2113] = 8'h08;	ram[2114] = 8'h23;	ram[2115] = 8'h34;
	ram[2116] = 8'hca;	ram[2117] = 8'ha4;	ram[2118] = 8'h08;	ram[2119] = 8'hcd;
	ram[2120] = 8'hd6;	ram[2121] = 8'h08;	ram[2122] = 8'hc3;	ram[2123] = 8'h7e;
	ram[2124] = 8'h08;	ram[2125] = 8'haf;	ram[2126] = 8'h90;	ram[2127] = 8'h47;
	ram[2128] = 8'h7e;	ram[2129] = 8'h9b;	ram[2130] = 8'h5f;	ram[2131] = 8'h23;
	ram[2132] = 8'h7e;	ram[2133] = 8'h9a;	ram[2134] = 8'h57;	ram[2135] = 8'h23;
	ram[2136] = 8'h7e;	ram[2137] = 8'h99;	ram[2138] = 8'h4f;	ram[2139] = 8'hdc;
	ram[2140] = 8'hb5;	ram[2141] = 8'h08;	ram[2142] = 8'h26;	ram[2143] = 8'h00;
	ram[2144] = 8'h79;	ram[2145] = 8'hb7;	ram[2146] = 8'hfa;	ram[2147] = 8'h7e;
	ram[2148] = 8'h08;	ram[2149] = 8'hfe;	ram[2150] = 8'he0;	ram[2151] = 8'hca;
	ram[2152] = 8'hbe;	ram[2153] = 8'h09;	ram[2154] = 8'h25;	ram[2155] = 8'h78;
	ram[2156] = 8'h87;	ram[2157] = 8'h47;	ram[2158] = 8'hcd;	ram[2159] = 8'h90;
	ram[2160] = 8'h08;	ram[2161] = 8'h7c;	ram[2162] = 8'hf2;	ram[2163] = 8'h65;
	ram[2164] = 8'h08;	ram[2165] = 8'h21;	ram[2166] = 8'h72;	ram[2167] = 8'h01;
	ram[2168] = 8'h86;	ram[2169] = 8'h77;	ram[2170] = 8'hd2;	ram[2171] = 8'hbe;
	ram[2172] = 8'h09;	ram[2173] = 8'hc8;	ram[2174] = 8'h78;	ram[2175] = 8'h21;
	ram[2176] = 8'h72;	ram[2177] = 8'h01;	ram[2178] = 8'hb7;	ram[2179] = 8'hfc;
	ram[2180] = 8'h9a;	ram[2181] = 8'h08;	ram[2182] = 8'h46;	ram[2183] = 8'h23;
	ram[2184] = 8'h7e;	ram[2185] = 8'he6;	ram[2186] = 8'h80;	ram[2187] = 8'ha9;
	ram[2188] = 8'h4f;	ram[2189] = 8'hc3;	ram[2190] = 8'h12;	ram[2191] = 8'h0a;
	ram[2192] = 8'h7b;	ram[2193] = 8'h17;	ram[2194] = 8'h5f;	ram[2195] = 8'h7a;
	ram[2196] = 8'h17;	ram[2197] = 8'h57;	ram[2198] = 8'h79;	ram[2199] = 8'h8f;
	ram[2200] = 8'h4f;	ram[2201] = 8'hc9;	ram[2202] = 8'h1c;	ram[2203] = 8'hc0;
	ram[2204] = 8'h14;	ram[2205] = 8'hc0;	ram[2206] = 8'h0c;	ram[2207] = 8'hc0;
	ram[2208] = 8'h0e;	ram[2209] = 8'h80;	ram[2210] = 8'h34;	ram[2211] = 8'hc0;
	ram[2212] = 8'h1e;	ram[2213] = 8'h0a;	ram[2214] = 8'hc3;	ram[2215] = 8'hd5;
	ram[2216] = 8'h01;	ram[2217] = 8'h7e;	ram[2218] = 8'h83;	ram[2219] = 8'h5f;
	ram[2220] = 8'h23;	ram[2221] = 8'h7e;	ram[2222] = 8'h8a;	ram[2223] = 8'h57;
	ram[2224] = 8'h23;	ram[2225] = 8'h7e;	ram[2226] = 8'h89;	ram[2227] = 8'h4f;
	ram[2228] = 8'hc9;	ram[2229] = 8'h21;	ram[2230] = 8'h73;	ram[2231] = 8'h01;
	ram[2232] = 8'h7e;	ram[2233] = 8'h2f;	ram[2234] = 8'h77;	ram[2235] = 8'haf;
	ram[2236] = 8'h6f;	ram[2237] = 8'h90;	ram[2238] = 8'h47;	ram[2239] = 8'h7d;
	ram[2240] = 8'h9b;	ram[2241] = 8'h5f;	ram[2242] = 8'h7d;	ram[2243] = 8'h9a;
	ram[2244] = 8'h57;	ram[2245] = 8'h7d;	ram[2246] = 8'h99;	ram[2247] = 8'h4f;
	ram[2248] = 8'hc9;	ram[2249] = 8'h06;	ram[2250] = 8'h00;	ram[2251] = 8'h3c;
	ram[2252] = 8'h6f;	ram[2253] = 8'haf;	ram[2254] = 8'h2d;	ram[2255] = 8'hc8;
	ram[2256] = 8'hcd;	ram[2257] = 8'hd6;	ram[2258] = 8'h08;	ram[2259] = 8'hc3;
	ram[2260] = 8'hcd;	ram[2261] = 8'h08;	ram[2262] = 8'h79;	ram[2263] = 8'h1f;
	ram[2264] = 8'h4f;	ram[2265] = 8'h7a;	ram[2266] = 8'h1f;	ram[2267] = 8'h57;
	ram[2268] = 8'h7b;	ram[2269] = 8'h1f;	ram[2270] = 8'h5f;	ram[2271] = 8'h78;
	ram[2272] = 8'h1f;	ram[2273] = 8'h47;	ram[2274] = 8'hc9;	ram[2275] = 8'hc1;
	ram[2276] = 8'hd1;	ram[2277] = 8'hef;	ram[2278] = 8'hc8;	ram[2279] = 8'h2e;
	ram[2280] = 8'h00;	ram[2281] = 8'hcd;	ram[2282] = 8'h9b;	ram[2283] = 8'h09;
	ram[2284] = 8'h79;	ram[2285] = 8'h32;	ram[2286] = 8'h17;	ram[2287] = 8'h09;
	ram[2288] = 8'heb;	ram[2289] = 8'h22;	ram[2290] = 8'h12;	ram[2291] = 8'h09;
	ram[2292] = 8'h01;	ram[2293] = 8'h00;	ram[2294] = 8'h00;	ram[2295] = 8'h50;
	ram[2296] = 8'h58;	ram[2297] = 8'h21;	ram[2298] = 8'h5e;	ram[2299] = 8'h08;
	ram[2300] = 8'he5;	ram[2301] = 8'h21;	ram[2302] = 8'h05;	ram[2303] = 8'h09;
	ram[2304] = 8'he5;	ram[2305] = 8'he5;	ram[2306] = 8'h21;	ram[2307] = 8'h6f;
	ram[2308] = 8'h01;	ram[2309] = 8'h7e;	ram[2310] = 8'h23;	ram[2311] = 8'he5;
	ram[2312] = 8'h2e;	ram[2313] = 8'h08;	ram[2314] = 8'h1f;	ram[2315] = 8'h67;
	ram[2316] = 8'h79;	ram[2317] = 8'hd2;	ram[2318] = 8'h19;	ram[2319] = 8'h09;
	ram[2320] = 8'he5;	ram[2321] = 8'h21;	ram[2322] = 8'h00;	ram[2323] = 8'h00;
	ram[2324] = 8'h19;	ram[2325] = 8'hd1;	ram[2326] = 8'hce;	ram[2327] = 8'h00;
	ram[2328] = 8'heb;	ram[2329] = 8'hcd;	ram[2330] = 8'hd7;	ram[2331] = 8'h08;
	ram[2332] = 8'h2d;	ram[2333] = 8'h7c;	ram[2334] = 8'hc2;	ram[2335] = 8'h0a;
	ram[2336] = 8'h09;	ram[2337] = 8'he1;	ram[2338] = 8'hc9;	ram[2339] = 8'hcd;
	ram[2340] = 8'h02;	ram[2341] = 8'h0a;	ram[2342] = 8'h01;	ram[2343] = 8'h20;
	ram[2344] = 8'h84;	ram[2345] = 8'h11;	ram[2346] = 8'h00;	ram[2347] = 8'h00;
	ram[2348] = 8'hcd;	ram[2349] = 8'h12;	ram[2350] = 8'h0a;	ram[2351] = 8'hc1;
	ram[2352] = 8'hd1;	ram[2353] = 8'hef;	ram[2354] = 8'hca;	ram[2355] = 8'hd3;
	ram[2356] = 8'h01;	ram[2357] = 8'h2e;	ram[2358] = 8'hff;	ram[2359] = 8'hcd;
	ram[2360] = 8'h9b;	ram[2361] = 8'h09;	ram[2362] = 8'h34;	ram[2363] = 8'h34;
	ram[2364] = 8'h2b;	ram[2365] = 8'h7e;	ram[2366] = 8'h32;	ram[2367] = 8'h60;
	ram[2368] = 8'h09;	ram[2369] = 8'h2b;	ram[2370] = 8'h7e;	ram[2371] = 8'h32;
	ram[2372] = 8'h5c;	ram[2373] = 8'h09;	ram[2374] = 8'h2b;	ram[2375] = 8'h7e;
	ram[2376] = 8'h32;	ram[2377] = 8'h58;	ram[2378] = 8'h09;	ram[2379] = 8'h41;
	ram[2380] = 8'heb;	ram[2381] = 8'haf;	ram[2382] = 8'h4f;	ram[2383] = 8'h57;
	ram[2384] = 8'h5f;	ram[2385] = 8'h32;	ram[2386] = 8'h63;	ram[2387] = 8'h09;
	ram[2388] = 8'he5;	ram[2389] = 8'hc5;	ram[2390] = 8'h7d;	ram[2391] = 8'hd6;
	ram[2392] = 8'h00;	ram[2393] = 8'h6f;	ram[2394] = 8'h7c;	ram[2395] = 8'hde;
	ram[2396] = 8'h00;	ram[2397] = 8'h67;	ram[2398] = 8'h78;	ram[2399] = 8'hde;
	ram[2400] = 8'h00;	ram[2401] = 8'h47;	ram[2402] = 8'h3e;	ram[2403] = 8'h00;
	ram[2404] = 8'hde;	ram[2405] = 8'h00;	ram[2406] = 8'h3f;	ram[2407] = 8'hd2;
	ram[2408] = 8'h71;	ram[2409] = 8'h09;	ram[2410] = 8'h32;	ram[2411] = 8'h63;
	ram[2412] = 8'h09;	ram[2413] = 8'hf1;	ram[2414] = 8'hf1;	ram[2415] = 8'h37;
	ram[2416] = 8'hd2;	ram[2417] = 8'hc1;	ram[2418] = 8'he1;	ram[2419] = 8'h79;
	ram[2420] = 8'h3c;	ram[2421] = 8'h3d;	ram[2422] = 8'h1f;	ram[2423] = 8'hfa;
	ram[2424] = 8'h7f;	ram[2425] = 8'h08;	ram[2426] = 8'h17;	ram[2427] = 8'hcd;
	ram[2428] = 8'h90;	ram[2429] = 8'h08;	ram[2430] = 8'h29;	ram[2431] = 8'h78;
	ram[2432] = 8'h17;	ram[2433] = 8'h47;	ram[2434] = 8'h3a;	ram[2435] = 8'h63;
	ram[2436] = 8'h09;	ram[2437] = 8'h17;	ram[2438] = 8'h32;	ram[2439] = 8'h63;
	ram[2440] = 8'h09;	ram[2441] = 8'h79;	ram[2442] = 8'hb2;	ram[2443] = 8'hb3;
	ram[2444] = 8'hc2;	ram[2445] = 8'h54;	ram[2446] = 8'h09;	ram[2447] = 8'he5;
	ram[2448] = 8'h21;	ram[2449] = 8'h72;	ram[2450] = 8'h01;	ram[2451] = 8'h35;
	ram[2452] = 8'he1;	ram[2453] = 8'hc2;	ram[2454] = 8'h54;	ram[2455] = 8'h09;
	ram[2456] = 8'hc3;	ram[2457] = 8'ha4;	ram[2458] = 8'h08;	ram[2459] = 8'h78;
	ram[2460] = 8'hb7;	ram[2461] = 8'hca;	ram[2462] = 8'hba;	ram[2463] = 8'h09;
	ram[2464] = 8'h7d;	ram[2465] = 8'h21;	ram[2466] = 8'h72;	ram[2467] = 8'h01;
	ram[2468] = 8'hae;	ram[2469] = 8'h80;	ram[2470] = 8'h47;	ram[2471] = 8'h1f;
	ram[2472] = 8'ha8;	ram[2473] = 8'h78;	ram[2474] = 8'hf2;	ram[2475] = 8'hb9;
	ram[2476] = 8'h09;	ram[2477] = 8'hc6;	ram[2478] = 8'h80;	ram[2479] = 8'h77;
	ram[2480] = 8'hca;	ram[2481] = 8'h21;	ram[2482] = 8'h09;	ram[2483] = 8'hcd;
	ram[2484] = 8'h37;	ram[2485] = 8'h0a;	ram[2486] = 8'h77;	ram[2487] = 8'h2b;
	ram[2488] = 8'hc9;	ram[2489] = 8'hb7;	ram[2490] = 8'he1;	ram[2491] = 8'hfa;
	ram[2492] = 8'ha4;	ram[2493] = 8'h08;	ram[2494] = 8'haf;	ram[2495] = 8'h32;
	ram[2496] = 8'h72;	ram[2497] = 8'h01;	ram[2498] = 8'hc9;	ram[2499] = 8'hcd;
	ram[2500] = 8'h1d;	ram[2501] = 8'h0a;	ram[2502] = 8'h78;	ram[2503] = 8'hb7;
	ram[2504] = 8'hc8;	ram[2505] = 8'hc6;	ram[2506] = 8'h02;	ram[2507] = 8'hda;
	ram[2508] = 8'ha4;	ram[2509] = 8'h08;	ram[2510] = 8'h47;	ram[2511] = 8'hcd;
	ram[2512] = 8'h12;	ram[2513] = 8'h08;	ram[2514] = 8'h21;	ram[2515] = 8'h72;
	ram[2516] = 8'h01;	ram[2517] = 8'h34;	ram[2518] = 8'hc0;	ram[2519] = 8'hc3;
	ram[2520] = 8'ha4;	ram[2521] = 8'h08;	ram[2522] = 8'h3a;	ram[2523] = 8'h71;
	ram[2524] = 8'h01;	ram[2525] = 8'hfe;	ram[2526] = 8'h2f;	ram[2527] = 8'h17;
	ram[2528] = 8'h9f;	ram[2529] = 8'hc0;	ram[2530] = 8'h3c;	ram[2531] = 8'hc9;
	ram[2532] = 8'hef;	ram[2533] = 8'h06;	ram[2534] = 8'h88;	ram[2535] = 8'h11;
	ram[2536] = 8'h00;	ram[2537] = 8'h00;	ram[2538] = 8'h21;	ram[2539] = 8'h72;
	ram[2540] = 8'h01;	ram[2541] = 8'h4f;	ram[2542] = 8'h70;	ram[2543] = 8'h06;
	ram[2544] = 8'h00;	ram[2545] = 8'h23;	ram[2546] = 8'h36;	ram[2547] = 8'h80;
	ram[2548] = 8'h17;	ram[2549] = 8'hc3;	ram[2550] = 8'h5b;	ram[2551] = 8'h08;
	ram[2552] = 8'hef;	ram[2553] = 8'hf0;	ram[2554] = 8'h21;	ram[2555] = 8'h71;
	ram[2556] = 8'h01;	ram[2557] = 8'h7e;	ram[2558] = 8'hee;	ram[2559] = 8'h80;
	ram[2560] = 8'h77;	ram[2561] = 8'hc9;	ram[2562] = 8'heb;	ram[2563] = 8'h2a;
	ram[2564] = 8'h6f;	ram[2565] = 8'h01;	ram[2566] = 8'he3;	ram[2567] = 8'he5;
	ram[2568] = 8'h2a;	ram[2569] = 8'h71;	ram[2570] = 8'h01;	ram[2571] = 8'he3;
	ram[2572] = 8'he5;	ram[2573] = 8'heb;	ram[2574] = 8'hc9;	ram[2575] = 8'hcd;
	ram[2576] = 8'h20;	ram[2577] = 8'h0a;	ram[2578] = 8'heb;	ram[2579] = 8'h22;
	ram[2580] = 8'h6f;	ram[2581] = 8'h01;	ram[2582] = 8'h60;	ram[2583] = 8'h69;
	ram[2584] = 8'h22;	ram[2585] = 8'h71;	ram[2586] = 8'h01;	ram[2587] = 8'heb;
	ram[2588] = 8'hc9;	ram[2589] = 8'h21;	ram[2590] = 8'h6f;	ram[2591] = 8'h01;
	ram[2592] = 8'h5e;	ram[2593] = 8'h23;	ram[2594] = 8'h56;	ram[2595] = 8'h23;
	ram[2596] = 8'h4e;	ram[2597] = 8'h23;	ram[2598] = 8'h46;	ram[2599] = 8'h23;
	ram[2600] = 8'hc9;	ram[2601] = 8'h11;	ram[2602] = 8'h6f;	ram[2603] = 8'h01;
	ram[2604] = 8'h06;	ram[2605] = 8'h04;	ram[2606] = 8'h1a;	ram[2607] = 8'h77;
	ram[2608] = 8'h13;	ram[2609] = 8'h23;	ram[2610] = 8'h05;	ram[2611] = 8'hc2;
	ram[2612] = 8'h2e;	ram[2613] = 8'h0a;	ram[2614] = 8'hc9;	ram[2615] = 8'h21;
	ram[2616] = 8'h71;	ram[2617] = 8'h01;	ram[2618] = 8'h7e;	ram[2619] = 8'h07;
	ram[2620] = 8'h37;	ram[2621] = 8'h1f;	ram[2622] = 8'h77;	ram[2623] = 8'h3f;
	ram[2624] = 8'h1f;	ram[2625] = 8'h23;	ram[2626] = 8'h23;	ram[2627] = 8'h77;
	ram[2628] = 8'h79;	ram[2629] = 8'h07;	ram[2630] = 8'h37;	ram[2631] = 8'h1f;
	ram[2632] = 8'h4f;	ram[2633] = 8'h1f;	ram[2634] = 8'hae;	ram[2635] = 8'hc9;
	ram[2636] = 8'h78;	ram[2637] = 8'hb7;	ram[2638] = 8'hca;	ram[2639] = 8'h28;
	ram[2640] = 8'h00;	ram[2641] = 8'h21;	ram[2642] = 8'hde;	ram[2643] = 8'h09;
	ram[2644] = 8'he5;	ram[2645] = 8'hef;	ram[2646] = 8'h79;	ram[2647] = 8'hc8;
	ram[2648] = 8'h21;	ram[2649] = 8'h71;	ram[2650] = 8'h01;	ram[2651] = 8'hae;
	ram[2652] = 8'h79;	ram[2653] = 8'hf8;	ram[2654] = 8'hcd;	ram[2655] = 8'h64;
	ram[2656] = 8'h0a;	ram[2657] = 8'h1f;	ram[2658] = 8'ha9;	ram[2659] = 8'hc9;
	ram[2660] = 8'h23;	ram[2661] = 8'h78;	ram[2662] = 8'hbe;	ram[2663] = 8'hc0;
	ram[2664] = 8'h2b;	ram[2665] = 8'h79;	ram[2666] = 8'hbe;	ram[2667] = 8'hc0;
	ram[2668] = 8'h2b;	ram[2669] = 8'h7a;	ram[2670] = 8'hbe;	ram[2671] = 8'hc0;
	ram[2672] = 8'h2b;	ram[2673] = 8'h7b;	ram[2674] = 8'h96;	ram[2675] = 8'hc0;
	ram[2676] = 8'he1;	ram[2677] = 8'he1;	ram[2678] = 8'hc9;	ram[2679] = 8'h47;
	ram[2680] = 8'h4f;	ram[2681] = 8'h57;	ram[2682] = 8'h5f;	ram[2683] = 8'hb7;
	ram[2684] = 8'hc8;	ram[2685] = 8'he5;	ram[2686] = 8'hcd;	ram[2687] = 8'h1d;
	ram[2688] = 8'h0a;	ram[2689] = 8'hcd;	ram[2690] = 8'h37;	ram[2691] = 8'h0a;
	ram[2692] = 8'hae;	ram[2693] = 8'h67;	ram[2694] = 8'hfc;	ram[2695] = 8'h9b;
	ram[2696] = 8'h0a;	ram[2697] = 8'h3e;	ram[2698] = 8'h98;	ram[2699] = 8'h90;
	ram[2700] = 8'hcd;	ram[2701] = 8'hc9;	ram[2702] = 8'h08;	ram[2703] = 8'h7c;
	ram[2704] = 8'h17;	ram[2705] = 8'hdc;	ram[2706] = 8'h9a;	ram[2707] = 8'h08;
	ram[2708] = 8'h06;	ram[2709] = 8'h00;	ram[2710] = 8'hdc;	ram[2711] = 8'hb5;
	ram[2712] = 8'h08;	ram[2713] = 8'he1;	ram[2714] = 8'hc9;	ram[2715] = 8'h1b;
	ram[2716] = 8'h7a;	ram[2717] = 8'ha3;	ram[2718] = 8'h3c;	ram[2719] = 8'hc0;
	ram[2720] = 8'h0d;	ram[2721] = 8'hc9;	ram[2722] = 8'h21;	ram[2723] = 8'h72;
	ram[2724] = 8'h01;	ram[2725] = 8'h7e;	ram[2726] = 8'hfe;	ram[2727] = 8'h98;
	ram[2728] = 8'hd0;	ram[2729] = 8'hcd;	ram[2730] = 8'h77;	ram[2731] = 8'h0a;
	ram[2732] = 8'h36;	ram[2733] = 8'h98;	ram[2734] = 8'h79;	ram[2735] = 8'h17;
	ram[2736] = 8'hc3;	ram[2737] = 8'h5b;	ram[2738] = 8'h08;	ram[2739] = 8'h2b;
	ram[2740] = 8'hcd;	ram[2741] = 8'hbe;	ram[2742] = 8'h09;	ram[2743] = 8'h47;
	ram[2744] = 8'h57;	ram[2745] = 8'h5f;	ram[2746] = 8'h2f;	ram[2747] = 8'h4f;
	ram[2748] = 8'hd7;	ram[2749] = 8'hda;	ram[2750] = 8'h04;	ram[2751] = 8'h0b;
	ram[2752] = 8'hfe;	ram[2753] = 8'h2e;	ram[2754] = 8'hca;	ram[2755] = 8'he4;
	ram[2756] = 8'h0a;	ram[2757] = 8'hfe;	ram[2758] = 8'h45;	ram[2759] = 8'hc2;
	ram[2760] = 8'he8;	ram[2761] = 8'h0a;	ram[2762] = 8'hd7;	ram[2763] = 8'h15;
	ram[2764] = 8'hfe;	ram[2765] = 8'h99;	ram[2766] = 8'hca;	ram[2767] = 8'hd8;
	ram[2768] = 8'h0a;	ram[2769] = 8'h14;	ram[2770] = 8'hfe;	ram[2771] = 8'h98;
	ram[2772] = 8'hca;	ram[2773] = 8'hd8;	ram[2774] = 8'h0a;	ram[2775] = 8'h2b;
	ram[2776] = 8'hd7;	ram[2777] = 8'hda;	ram[2778] = 8'h23;	ram[2779] = 8'h0b;
	ram[2780] = 8'h14;	ram[2781] = 8'hc2;	ram[2782] = 8'he8;	ram[2783] = 8'h0a;
	ram[2784] = 8'haf;	ram[2785] = 8'h93;	ram[2786] = 8'h5f;	ram[2787] = 8'h0c;
	ram[2788] = 8'h0c;	ram[2789] = 8'hca;	ram[2790] = 8'hbc;	ram[2791] = 8'h0a;
	ram[2792] = 8'he5;	ram[2793] = 8'h7b;	ram[2794] = 8'h90;	ram[2795] = 8'hf4;
	ram[2796] = 8'hfc;	ram[2797] = 8'h0a;	ram[2798] = 8'hf2;	ram[2799] = 8'hf7;
	ram[2800] = 8'h0a;	ram[2801] = 8'hf5;	ram[2802] = 8'hcd;	ram[2803] = 8'h23;
	ram[2804] = 8'h09;	ram[2805] = 8'hf1;	ram[2806] = 8'h3c;	ram[2807] = 8'hc2;
	ram[2808] = 8'heb;	ram[2809] = 8'h0a;	ram[2810] = 8'he1;	ram[2811] = 8'hc9;
	ram[2812] = 8'hc8;	ram[2813] = 8'hf5;	ram[2814] = 8'hcd;	ram[2815] = 8'hc3;
	ram[2816] = 8'h09;	ram[2817] = 8'hf1;	ram[2818] = 8'h3d;	ram[2819] = 8'hc9;
	ram[2820] = 8'hd5;	ram[2821] = 8'h57;	ram[2822] = 8'h78;	ram[2823] = 8'h89;
	ram[2824] = 8'h47;	ram[2825] = 8'hc5;	ram[2826] = 8'he5;	ram[2827] = 8'hd5;
	ram[2828] = 8'hcd;	ram[2829] = 8'hc3;	ram[2830] = 8'h09;	ram[2831] = 8'hf1;
	ram[2832] = 8'hd6;	ram[2833] = 8'h30;	ram[2834] = 8'hcd;	ram[2835] = 8'h02;
	ram[2836] = 8'h0a;	ram[2837] = 8'hcd;	ram[2838] = 8'he5;	ram[2839] = 8'h09;
	ram[2840] = 8'hc1;	ram[2841] = 8'hd1;	ram[2842] = 8'hcd;	ram[2843] = 8'h12;
	ram[2844] = 8'h08;	ram[2845] = 8'he1;	ram[2846] = 8'hc1;	ram[2847] = 8'hd1;
	ram[2848] = 8'hc3;	ram[2849] = 8'hbc;	ram[2850] = 8'h0a;	ram[2851] = 8'h7b;
	ram[2852] = 8'h07;	ram[2853] = 8'h07;	ram[2854] = 8'h83;	ram[2855] = 8'h07;
	ram[2856] = 8'h86;	ram[2857] = 8'hd6;	ram[2858] = 8'h30;	ram[2859] = 8'h5f;
	ram[2860] = 8'hc3;	ram[2861] = 8'hd8;	ram[2862] = 8'h0a;	ram[2863] = 8'he5;
	ram[2864] = 8'h21;	ram[2865] = 8'h88;	ram[2866] = 8'h01;	ram[2867] = 8'hcd;
	ram[2868] = 8'ha3;	ram[2869] = 8'h05;	ram[2870] = 8'he1;	ram[2871] = 8'heb;
	ram[2872] = 8'haf;	ram[2873] = 8'h06;	ram[2874] = 8'h98;	ram[2875] = 8'hcd;
	ram[2876] = 8'hea;	ram[2877] = 8'h09;	ram[2878] = 8'h21;	ram[2879] = 8'ha2;
	ram[2880] = 8'h05;	ram[2881] = 8'he5;	ram[2882] = 8'h21;	ram[2883] = 8'h74;
	ram[2884] = 8'h01;	ram[2885] = 8'he5;	ram[2886] = 8'hef;	ram[2887] = 8'h36;
	ram[2888] = 8'h20;	ram[2889] = 8'hf2;	ram[2890] = 8'h4e;	ram[2891] = 8'h0b;
	ram[2892] = 8'h36;	ram[2893] = 8'h2d;	ram[2894] = 8'h23;	ram[2895] = 8'h36;
	ram[2896] = 8'h30;	ram[2897] = 8'hca;	ram[2898] = 8'hf7;	ram[2899] = 8'h0b;
	ram[2900] = 8'he5;	ram[2901] = 8'hfc;	ram[2902] = 8'hfa;	ram[2903] = 8'h09;
	ram[2904] = 8'haf;	ram[2905] = 8'hf5;	ram[2906] = 8'hcd;	ram[2907] = 8'hfd;
	ram[2908] = 8'h0b;	ram[2909] = 8'h01;	ram[2910] = 8'h43;	ram[2911] = 8'h91;
	ram[2912] = 8'h11;	ram[2913] = 8'hf8;	ram[2914] = 8'h4f;	ram[2915] = 8'hcd;
	ram[2916] = 8'h4c;	ram[2917] = 8'h0a;	ram[2918] = 8'he2;	ram[2919] = 8'h7a;
	ram[2920] = 8'h0b;	ram[2921] = 8'hf1;	ram[2922] = 8'hcd;	ram[2923] = 8'hfd;
	ram[2924] = 8'h0a;	ram[2925] = 8'hf5;	ram[2926] = 8'hc3;	ram[2927] = 8'h5d;
	ram[2928] = 8'h0b;	ram[2929] = 8'hcd;	ram[2930] = 8'h23;	ram[2931] = 8'h09;
	ram[2932] = 8'hf1;	ram[2933] = 8'h3c;	ram[2934] = 8'hf5;	ram[2935] = 8'hcd;
	ram[2936] = 8'hfd;	ram[2937] = 8'h0b;	ram[2938] = 8'hcd;	ram[2939] = 8'h01;
	ram[2940] = 8'h08;	ram[2941] = 8'h3c;	ram[2942] = 8'hcd;	ram[2943] = 8'h77;
	ram[2944] = 8'h0a;	ram[2945] = 8'hcd;	ram[2946] = 8'h12;	ram[2947] = 8'h0a;
	ram[2948] = 8'h01;	ram[2949] = 8'h06;	ram[2950] = 8'h02;	ram[2951] = 8'hf1;
	ram[2952] = 8'h81;	ram[2953] = 8'hfa;	ram[2954] = 8'h95;	ram[2955] = 8'h0b;
	ram[2956] = 8'hfe;	ram[2957] = 8'h07;	ram[2958] = 8'hd2;	ram[2959] = 8'h95;
	ram[2960] = 8'h0b;	ram[2961] = 8'h3c;	ram[2962] = 8'h47;	ram[2963] = 8'h3e;
	ram[2964] = 8'h01;	ram[2965] = 8'h3d;	ram[2966] = 8'he1;	ram[2967] = 8'hf5;
	ram[2968] = 8'h11;	ram[2969] = 8'h0f;	ram[2970] = 8'h0c;	ram[2971] = 8'h05;
	ram[2972] = 8'h36;	ram[2973] = 8'h2e;	ram[2974] = 8'hcc;	ram[2975] = 8'h27;
	ram[2976] = 8'h0a;	ram[2977] = 8'hc5;	ram[2978] = 8'he5;	ram[2979] = 8'hd5;
	ram[2980] = 8'hcd;	ram[2981] = 8'h1d;	ram[2982] = 8'h0a;	ram[2983] = 8'he1;
	ram[2984] = 8'h06;	ram[2985] = 8'h2f;	ram[2986] = 8'h04;	ram[2987] = 8'h7b;
	ram[2988] = 8'h96;	ram[2989] = 8'h5f;	ram[2990] = 8'h23;	ram[2991] = 8'h7a;
	ram[2992] = 8'h9e;	ram[2993] = 8'h57;	ram[2994] = 8'h23;	ram[2995] = 8'h79;
	ram[2996] = 8'h9e;	ram[2997] = 8'h4f;	ram[2998] = 8'h2b;	ram[2999] = 8'h2b;
	ram[3000] = 8'hd2;	ram[3001] = 8'haa;	ram[3002] = 8'h0b;	ram[3003] = 8'hcd;
	ram[3004] = 8'ha9;	ram[3005] = 8'h08;	ram[3006] = 8'h23;	ram[3007] = 8'hcd;
	ram[3008] = 8'h12;	ram[3009] = 8'h0a;	ram[3010] = 8'heb;	ram[3011] = 8'he1;
	ram[3012] = 8'h70;	ram[3013] = 8'h23;	ram[3014] = 8'hc1;	ram[3015] = 8'h0d;
	ram[3016] = 8'hc2;	ram[3017] = 8'h9b;	ram[3018] = 8'h0b;	ram[3019] = 8'h05;
	ram[3020] = 8'hca;	ram[3021] = 8'hdb;	ram[3022] = 8'h0b;	ram[3023] = 8'h2b;
	ram[3024] = 8'h7e;	ram[3025] = 8'hfe;	ram[3026] = 8'h30;	ram[3027] = 8'hca;
	ram[3028] = 8'hcf;	ram[3029] = 8'h0b;	ram[3030] = 8'hfe;	ram[3031] = 8'h2e;
	ram[3032] = 8'hc4;	ram[3033] = 8'h27;	ram[3034] = 8'h0a;	ram[3035] = 8'hf1;
	ram[3036] = 8'hca;	ram[3037] = 8'hfa;	ram[3038] = 8'h0b;	ram[3039] = 8'h36;
	ram[3040] = 8'h45;	ram[3041] = 8'h23;	ram[3042] = 8'h36;	ram[3043] = 8'h2b;
	ram[3044] = 8'hf2;	ram[3045] = 8'heb;	ram[3046] = 8'h0b;	ram[3047] = 8'h36;
	ram[3048] = 8'h2d;	ram[3049] = 8'h2f;	ram[3050] = 8'h3c;	ram[3051] = 8'h06;
	ram[3052] = 8'h2f;	ram[3053] = 8'h04;	ram[3054] = 8'hd6;	ram[3055] = 8'h0a;
	ram[3056] = 8'hd2;	ram[3057] = 8'hed;	ram[3058] = 8'h0b;	ram[3059] = 8'hc6;
	ram[3060] = 8'h3a;	ram[3061] = 8'h23;	ram[3062] = 8'h70;	ram[3063] = 8'h23;
	ram[3064] = 8'h77;	ram[3065] = 8'h23;	ram[3066] = 8'h71;	ram[3067] = 8'he1;
	ram[3068] = 8'hc9;	ram[3069] = 8'h01;	ram[3070] = 8'h74;	ram[3071] = 8'h94;
	ram[3072] = 8'h11;	ram[3073] = 8'hf7;	ram[3074] = 8'h23;	ram[3075] = 8'hcd;
	ram[3076] = 8'h4c;	ram[3077] = 8'h0a;	ram[3078] = 8'he1;	ram[3079] = 8'he2;
	ram[3080] = 8'h71;	ram[3081] = 8'h0b;	ram[3082] = 8'he9;	ram[3083] = 8'h00;
	ram[3084] = 8'h00;	ram[3085] = 8'h00;	ram[3086] = 8'h80;	ram[3087] = 8'ha0;
	ram[3088] = 8'h86;	ram[3089] = 8'h01;	ram[3090] = 8'h10;	ram[3091] = 8'h27;
	ram[3092] = 8'h00;	ram[3093] = 8'he8;	ram[3094] = 8'h03;	ram[3095] = 8'h00;
	ram[3096] = 8'h64;	ram[3097] = 8'h00;	ram[3098] = 8'h00;	ram[3099] = 8'h0a;
	ram[3100] = 8'h00;	ram[3101] = 8'h00;	ram[3102] = 8'h01;	ram[3103] = 8'h00;
	ram[3104] = 8'h00;	ram[3105] = 8'hef;	ram[3106] = 8'hfa;	ram[3107] = 8'h98;
	ram[3108] = 8'h04;	ram[3109] = 8'hc8;	ram[3110] = 8'h21;	ram[3111] = 8'h72;
	ram[3112] = 8'h01;	ram[3113] = 8'h7e;	ram[3114] = 8'h1f;	ram[3115] = 8'hf5;
	ram[3116] = 8'he5;	ram[3117] = 8'h3e;	ram[3118] = 8'h40;	ram[3119] = 8'h17;
	ram[3120] = 8'h77;	ram[3121] = 8'h21;	ram[3122] = 8'h74;	ram[3123] = 8'h01;
	ram[3124] = 8'hcd;	ram[3125] = 8'h29;	ram[3126] = 8'h0a;	ram[3127] = 8'h3e;
	ram[3128] = 8'h04;	ram[3129] = 8'hf5;	ram[3130] = 8'hcd;	ram[3131] = 8'h02;
	ram[3132] = 8'h0a;	ram[3133] = 8'h21;	ram[3134] = 8'h74;	ram[3135] = 8'h01;
	ram[3136] = 8'hcd;	ram[3137] = 8'h20;	ram[3138] = 8'h0a;	ram[3139] = 8'hcd;
	ram[3140] = 8'h31;	ram[3141] = 8'h09;	ram[3142] = 8'hc1;	ram[3143] = 8'hd1;
	ram[3144] = 8'hcd;	ram[3145] = 8'h12;	ram[3146] = 8'h08;	ram[3147] = 8'h01;
	ram[3148] = 8'h00;	ram[3149] = 8'h80;	ram[3150] = 8'h51;	ram[3151] = 8'h59;
	ram[3152] = 8'hcd;	ram[3153] = 8'he5;	ram[3154] = 8'h08;	ram[3155] = 8'hf1;
	ram[3156] = 8'h3d;	ram[3157] = 8'hc2;	ram[3158] = 8'h39;	ram[3159] = 8'h0c;
	ram[3160] = 8'he1;	ram[3161] = 8'hf1;	ram[3162] = 8'hc6;	ram[3163] = 8'hc0;
	ram[3164] = 8'h86;	ram[3165] = 8'h77;	ram[3166] = 8'hc9;	ram[3167] = 8'hef;
	ram[3168] = 8'hfa;	ram[3169] = 8'h7c;	ram[3170] = 8'h0c;	ram[3171] = 8'h21;
	ram[3172] = 8'h91;	ram[3173] = 8'h0c;	ram[3174] = 8'hcd;	ram[3175] = 8'h0f;
	ram[3176] = 8'h0a;	ram[3177] = 8'hc8;	ram[3178] = 8'h01;	ram[3179] = 8'h35;
	ram[3180] = 8'h98;	ram[3181] = 8'h11;	ram[3182] = 8'h7a;	ram[3183] = 8'h44;
	ram[3184] = 8'hcd;	ram[3185] = 8'he5;	ram[3186] = 8'h08;	ram[3187] = 8'h01;
	ram[3188] = 8'h28;	ram[3189] = 8'h68;	ram[3190] = 8'h11;	ram[3191] = 8'h46;
	ram[3192] = 8'hb1;	ram[3193] = 8'hcd;	ram[3194] = 8'h12;	ram[3195] = 8'h08;
	ram[3196] = 8'hcd;	ram[3197] = 8'h1d;	ram[3198] = 8'h0a;	ram[3199] = 8'h7b;
	ram[3200] = 8'h59;	ram[3201] = 8'h4f;	ram[3202] = 8'h36;	ram[3203] = 8'h80;
	ram[3204] = 8'h2b;	ram[3205] = 8'h46;	ram[3206] = 8'h36;	ram[3207] = 8'h80;
	ram[3208] = 8'hcd;	ram[3209] = 8'h5e;	ram[3210] = 8'h08;	ram[3211] = 8'h21;
	ram[3212] = 8'h91;	ram[3213] = 8'h0c;	ram[3214] = 8'hc3;	ram[3215] = 8'h29;
	ram[3216] = 8'h0a;	ram[3217] = 8'h52;	ram[3218] = 8'hc7;	ram[3219] = 8'h4f;
	ram[3220] = 8'h80;	ram[3221] = 8'hcd;	ram[3222] = 8'h02;	ram[3223] = 8'h0a;
	ram[3224] = 8'h01;	ram[3225] = 8'h49;	ram[3226] = 8'h83;	ram[3227] = 8'h11;
	ram[3228] = 8'hdb;	ram[3229] = 8'h0f;	ram[3230] = 8'hcd;	ram[3231] = 8'h12;
	ram[3232] = 8'h0a;	ram[3233] = 8'hc1;	ram[3234] = 8'hd1;	ram[3235] = 8'hcd;
	ram[3236] = 8'h31;	ram[3237] = 8'h09;	ram[3238] = 8'hcd;	ram[3239] = 8'h02;
	ram[3240] = 8'h0a;	ram[3241] = 8'hcd;	ram[3242] = 8'ha2;	ram[3243] = 8'h0a;
	ram[3244] = 8'hc1;	ram[3245] = 8'hd1;	ram[3246] = 8'hcd;	ram[3247] = 8'h0c;
	ram[3248] = 8'h08;	ram[3249] = 8'h01;	ram[3250] = 8'h00;	ram[3251] = 8'h7f;
	ram[3252] = 8'h51;	ram[3253] = 8'h59;	ram[3254] = 8'hcd;	ram[3255] = 8'h0c;
	ram[3256] = 8'h08;	ram[3257] = 8'hef;	ram[3258] = 8'h37;	ram[3259] = 8'hf2;
	ram[3260] = 8'hc3;	ram[3261] = 8'h0c;	ram[3262] = 8'hcd;	ram[3263] = 8'h01;
	ram[3264] = 8'h08;	ram[3265] = 8'hef;	ram[3266] = 8'hb7;	ram[3267] = 8'hf5;
	ram[3268] = 8'hf4;	ram[3269] = 8'hfa;	ram[3270] = 8'h09;	ram[3271] = 8'h01;
	ram[3272] = 8'h00;	ram[3273] = 8'h7f;	ram[3274] = 8'h51;	ram[3275] = 8'h59;
	ram[3276] = 8'hcd;	ram[3277] = 8'h12;	ram[3278] = 8'h08;	ram[3279] = 8'hf1;
	ram[3280] = 8'hd4;	ram[3281] = 8'hfa;	ram[3282] = 8'h09;	ram[3283] = 8'hcd;
	ram[3284] = 8'h02;	ram[3285] = 8'h0a;	ram[3286] = 8'hcd;	ram[3287] = 8'h1d;
	ram[3288] = 8'h0a;	ram[3289] = 8'hcd;	ram[3290] = 8'he5;	ram[3291] = 8'h08;
	ram[3292] = 8'hcd;	ram[3293] = 8'h02;	ram[3294] = 8'h0a;	ram[3295] = 8'h21;
	ram[3296] = 8'h03;	ram[3297] = 8'h0d;	ram[3298] = 8'hcd;	ram[3299] = 8'h0f;
	ram[3300] = 8'h0a;	ram[3301] = 8'hc1;	ram[3302] = 8'hd1;	ram[3303] = 8'h3e;
	ram[3304] = 8'h04;	ram[3305] = 8'hf5;	ram[3306] = 8'hd5;	ram[3307] = 8'hc5;
	ram[3308] = 8'he5;	ram[3309] = 8'hcd;	ram[3310] = 8'he5;	ram[3311] = 8'h08;
	ram[3312] = 8'he1;	ram[3313] = 8'hcd;	ram[3314] = 8'h20;	ram[3315] = 8'h0a;
	ram[3316] = 8'he5;	ram[3317] = 8'hcd;	ram[3318] = 8'h12;	ram[3319] = 8'h08;
	ram[3320] = 8'he1;	ram[3321] = 8'hc1;	ram[3322] = 8'hd1;	ram[3323] = 8'hf1;
	ram[3324] = 8'h3d;	ram[3325] = 8'hc2;	ram[3326] = 8'he9;	ram[3327] = 8'h0c;
	ram[3328] = 8'hc3;	ram[3329] = 8'he3;	ram[3330] = 8'h08;	ram[3331] = 8'hba;
	ram[3332] = 8'hd7;	ram[3333] = 8'h1e;	ram[3334] = 8'h86;	ram[3335] = 8'h64;
	ram[3336] = 8'h26;	ram[3337] = 8'h99;	ram[3338] = 8'h87;	ram[3339] = 8'h58;
	ram[3340] = 8'h34;	ram[3341] = 8'h23;	ram[3342] = 8'h87;	ram[3343] = 8'he0;
	ram[3344] = 8'h5d;	ram[3345] = 8'ha5;	ram[3346] = 8'h86;	ram[3347] = 8'hda;
	ram[3348] = 8'h0f;	ram[3349] = 8'h49;	ram[3350] = 8'h83;	ram[3351] = 8'h00;
	ram[3352] = 8'h00;	ram[3353] = 8'h00;	ram[3354] = 8'h00;	ram[3355] = 8'h00;
	ram[3356] = 8'h00;	ram[3357] = 8'h00;	ram[3358] = 8'h00;	ram[3359] = 8'h00;
	ram[3360] = 8'h00;	ram[3361] = 8'h21;	ram[3362] = 8'h1a;	ram[3363] = 8'h0f;
	ram[3364] = 8'hf9;	ram[3365] = 8'h22;	ram[3366] = 8'h63;	ram[3367] = 8'h01;
	ram[3368] = 8'hdb;	ram[3369] = 8'h01;	ram[3370] = 8'h0e;	ram[3371] = 8'hff;
	ram[3372] = 8'h11;	ram[3373] = 8'h8e;	ram[3374] = 8'h0d;	ram[3375] = 8'hd5;
	ram[3376] = 8'h3a;	ram[3377] = 8'hff;	ram[3378] = 8'h0f;	ram[3379] = 8'h47;
	ram[3380] = 8'hdb;	ram[3381] = 8'hff;	ram[3382] = 8'h1f;	ram[3383] = 8'hda;
	ram[3384] = 8'h41;	ram[3385] = 8'h0d;	ram[3386] = 8'he6;	ram[3387] = 8'h0c;
	ram[3388] = 8'hca;	ram[3389] = 8'h42;	ram[3390] = 8'h0d;	ram[3391] = 8'h06;
	ram[3392] = 8'h10;	ram[3393] = 8'h78;	ram[3394] = 8'h32;	ram[3395] = 8'h8c;
	ram[3396] = 8'h0d;	ram[3397] = 8'hdb;	ram[3398] = 8'hff;	ram[3399] = 8'h17;
	ram[3400] = 8'h17;	ram[3401] = 8'h06;	ram[3402] = 8'h20;	ram[3403] = 8'h11;
	ram[3404] = 8'h02;	ram[3405] = 8'hca;	ram[3406] = 8'hd8;	ram[3407] = 8'h17;
	ram[3408] = 8'h43;	ram[3409] = 8'h1d;	ram[3410] = 8'hd8;	ram[3411] = 8'h17;
	ram[3412] = 8'hda;	ram[3413] = 8'h6f;	ram[3414] = 8'h0d;	ram[3415] = 8'h43;
	ram[3416] = 8'h11;	ram[3417] = 8'h80;	ram[3418] = 8'hc2;	ram[3419] = 8'h17;
	ram[3420] = 8'hd0;	ram[3421] = 8'h17;	ram[3422] = 8'h3e;	ram[3423] = 8'h03;
	ram[3424] = 8'hcd;	ram[3425] = 8'h8b;	ram[3426] = 8'h0d;	ram[3427] = 8'h3d;
	ram[3428] = 8'h8f;	ram[3429] = 8'h87;	ram[3430] = 8'h87;	ram[3431] = 8'h3c;
	ram[3432] = 8'hcd;	ram[3433] = 8'h8b;	ram[3434] = 8'h0d;	ram[3435] = 8'h37;
	ram[3436] = 8'hc3;	ram[3437] = 8'h4b;	ram[3438] = 8'h0d;	ram[3439] = 8'haf;
	ram[3440] = 8'hcd;	ram[3441] = 8'h8b;	ram[3442] = 8'h0d;	ram[3443] = 8'hcd;
	ram[3444] = 8'h87;	ram[3445] = 8'h0d;	ram[3446] = 8'hcd;	ram[3447] = 8'h87;
	ram[3448] = 8'h0d;	ram[3449] = 8'h4b;	ram[3450] = 8'h2f;	ram[3451] = 8'hcd;
	ram[3452] = 8'h87;	ram[3453] = 8'h0d;	ram[3454] = 8'h3e;	ram[3455] = 8'h04;
	ram[3456] = 8'h35;	ram[3457] = 8'hcd;	ram[3458] = 8'h8b;	ram[3459] = 8'h0d;
	ram[3460] = 8'h35;	ram[3461] = 8'h35;	ram[3462] = 8'h35;	ram[3463] = 8'h21;
	ram[3464] = 8'h8c;	ram[3465] = 8'h0d;	ram[3466] = 8'h34;	ram[3467] = 8'hd3;
	ram[3468] = 8'h10;	ram[3469] = 8'hc9;	ram[3470] = 8'h62;	ram[3471] = 8'h68;
	ram[3472] = 8'h22;	ram[3473] = 8'h85;	ram[3474] = 8'h03;	ram[3475] = 8'h7c;
	ram[3476] = 8'he6;	ram[3477] = 8'hc8;	ram[3478] = 8'h67;	ram[3479] = 8'h22;
	ram[3480] = 8'h76;	ram[3481] = 8'h04;	ram[3482] = 8'heb;	ram[3483] = 8'h22;
	ram[3484] = 8'h7a;	ram[3485] = 8'h03;	ram[3486] = 8'h3a;	ram[3487] = 8'h8c;
	ram[3488] = 8'h0d;	ram[3489] = 8'h32;	ram[3490] = 8'h83;	ram[3491] = 8'h03;
	ram[3492] = 8'h32;	ram[3493] = 8'h74;	ram[3494] = 8'h04;	ram[3495] = 8'h3c;
	ram[3496] = 8'h32;	ram[3497] = 8'h8a;	ram[3498] = 8'h03;	ram[3499] = 8'h81;
	ram[3500] = 8'h32;	ram[3501] = 8'h78;	ram[3502] = 8'h03;	ram[3503] = 8'h3c;
	ram[3504] = 8'h32;	ram[3505] = 8'h80;	ram[3506] = 8'h03;	ram[3507] = 8'h21;
	ram[3508] = 8'hff;	ram[3509] = 8'hff;	ram[3510] = 8'h22;	ram[3511] = 8'h61;
	ram[3512] = 8'h01;	ram[3513] = 8'hcd;	ram[3514] = 8'h8a;	ram[3515] = 8'h05;
	ram[3516] = 8'h21;	ram[3517] = 8'hf0;	ram[3518] = 8'h0e;	ram[3519] = 8'hcd;
	ram[3520] = 8'ha3;	ram[3521] = 8'h05;	ram[3522] = 8'hcd;	ram[3523] = 8'hc2;
	ram[3524] = 8'h02;	ram[3525] = 8'hd7;	ram[3526] = 8'hb7;	ram[3527] = 8'hc2;
	ram[3528] = 8'hde;	ram[3529] = 8'h0d;	ram[3530] = 8'h21;	ram[3531] = 8'hfc;
	ram[3532] = 8'h0e;	ram[3533] = 8'h23;	ram[3534] = 8'h3e;	ram[3535] = 8'h37;
	ram[3536] = 8'h77;	ram[3537] = 8'hbe;	ram[3538] = 8'hc2;	ram[3539] = 8'hea;
	ram[3540] = 8'h0d;	ram[3541] = 8'h3d;	ram[3542] = 8'h77;	ram[3543] = 8'hbe;
	ram[3544] = 8'hca;	ram[3545] = 8'hcd;	ram[3546] = 8'h0d;	ram[3547] = 8'hc3;
	ram[3548] = 8'hea;	ram[3549] = 8'h0d;	ram[3550] = 8'h21;	ram[3551] = 8'h13;
	ram[3552] = 8'h01;	ram[3553] = 8'hcd;	ram[3554] = 8'h9d;	ram[3555] = 8'h04;
	ram[3556] = 8'hb7;	ram[3557] = 8'hc2;	ram[3558] = 8'hd0;	ram[3559] = 8'h01;
	ram[3560] = 8'heb;	ram[3561] = 8'h2b;	ram[3562] = 8'h2b;	ram[3563] = 8'he5;
	ram[3564] = 8'h21;	ram[3565] = 8'hb4;	ram[3566] = 8'h0e;	ram[3567] = 8'hcd;
	ram[3568] = 8'ha3;	ram[3569] = 8'h05;	ram[3570] = 8'hcd;	ram[3571] = 8'hc2;
	ram[3572] = 8'h02;	ram[3573] = 8'hd7;	ram[3574] = 8'hb7;	ram[3575] = 8'hca;
	ram[3576] = 8'h1b;	ram[3577] = 8'h0e;	ram[3578] = 8'h21;	ram[3579] = 8'h13;
	ram[3580] = 8'h01;	ram[3581] = 8'hcd;	ram[3582] = 8'h9d;	ram[3583] = 8'h04;
	ram[3584] = 8'h7a;	ram[3585] = 8'hb7;	ram[3586] = 8'hc2;	ram[3587] = 8'hec;
	ram[3588] = 8'h0d;	ram[3589] = 8'h7b;	ram[3590] = 8'hfe;	ram[3591] = 8'h10;
	ram[3592] = 8'hda;	ram[3593] = 8'hec;	ram[3594] = 8'h0d;	ram[3595] = 8'h32;
	ram[3596] = 8'h6f;	ram[3597] = 8'h03;	ram[3598] = 8'hd6;	ram[3599] = 8'h0e;
	ram[3600] = 8'hd2;	ram[3601] = 8'h0e;	ram[3602] = 8'h0e;	ram[3603] = 8'hc6;
	ram[3604] = 8'h1c;	ram[3605] = 8'h2f;	ram[3606] = 8'h3c;	ram[3607] = 8'h83;
	ram[3608] = 8'h32;	ram[3609] = 8'hb7;	ram[3610] = 8'h05;	ram[3611] = 8'h21;
	ram[3612] = 8'h85;	ram[3613] = 8'h0e;	ram[3614] = 8'hf7;	ram[3615] = 8'h11;
	ram[3616] = 8'h99;	ram[3617] = 8'h0e;	ram[3618] = 8'he7;	ram[3619] = 8'hca;
	ram[3620] = 8'h32;	ram[3621] = 8'h0e;	ram[3622] = 8'hf7;	ram[3623] = 8'he3;
	ram[3624] = 8'hcd;	ram[3625] = 8'ha3;	ram[3626] = 8'h05;	ram[3627] = 8'hcd;
	ram[3628] = 8'hc2;	ram[3629] = 8'h02;	ram[3630] = 8'hd7;	ram[3631] = 8'he1;
	ram[3632] = 8'hfe;	ram[3633] = 8'h59;	ram[3634] = 8'hd1;	ram[3635] = 8'hca;
	ram[3636] = 8'h47;	ram[3637] = 8'h0e;	ram[3638] = 8'hfe;	ram[3639] = 8'h4e;
	ram[3640] = 8'hc2;	ram[3641] = 8'h1b;	ram[3642] = 8'h0e;	ram[3643] = 8'hf7;
	ram[3644] = 8'he3;	ram[3645] = 8'h11;	ram[3646] = 8'h98;	ram[3647] = 8'h04;
	ram[3648] = 8'h73;	ram[3649] = 8'h23;	ram[3650] = 8'h72;	ram[3651] = 8'he1;
	ram[3652] = 8'hc3;	ram[3653] = 8'h1e;	ram[3654] = 8'h0e;	ram[3655] = 8'heb;
	ram[3656] = 8'h36;	ram[3657] = 8'h00;	ram[3658] = 8'h23;	ram[3659] = 8'h22;
	ram[3660] = 8'h65;	ram[3661] = 8'h01;	ram[3662] = 8'he3;	ram[3663] = 8'h11;
	ram[3664] = 8'h1a;	ram[3665] = 8'h0f;	ram[3666] = 8'he7;	ram[3667] = 8'hda;
	ram[3668] = 8'hcd;	ram[3669] = 8'h01;	ram[3670] = 8'hd1;	ram[3671] = 8'hf9;
	ram[3672] = 8'h22;	ram[3673] = 8'h63;	ram[3674] = 8'h01;	ram[3675] = 8'heb;
	ram[3676] = 8'hcd;	ram[3677] = 8'hc3;	ram[3678] = 8'h01;	ram[3679] = 8'h7b;
	ram[3680] = 8'h95;	ram[3681] = 8'h6f;	ram[3682] = 8'h7a;	ram[3683] = 8'h9c;
	ram[3684] = 8'h67;	ram[3685] = 8'h01;	ram[3686] = 8'hf0;	ram[3687] = 8'hff;
	ram[3688] = 8'h09;	ram[3689] = 8'hcd;	ram[3690] = 8'h8a;	ram[3691] = 8'h05;
	ram[3692] = 8'hcd;	ram[3693] = 8'h37;	ram[3694] = 8'h0b;	ram[3695] = 8'h21;
	ram[3696] = 8'hc3;	ram[3697] = 8'h0e;	ram[3698] = 8'hcd;	ram[3699] = 8'ha3;
	ram[3700] = 8'h05;	ram[3701] = 8'h21;	ram[3702] = 8'ha3;	ram[3703] = 8'h05;
	ram[3704] = 8'h22;	ram[3705] = 8'hfd;	ram[3706] = 8'h01;	ram[3707] = 8'hcd;
	ram[3708] = 8'h96;	ram[3709] = 8'h02;	ram[3710] = 8'h21;	ram[3711] = 8'hf9;
	ram[3712] = 8'h01;	ram[3713] = 8'h22;	ram[3714] = 8'h02;	ram[3715] = 8'h00;
	ram[3716] = 8'he9;	ram[3717] = 8'h17;	ram[3718] = 8'h0d;	ram[3719] = 8'h99;
	ram[3720] = 8'h0e;	ram[3721] = 8'h49;	ram[3722] = 8'h00;	ram[3723] = 8'h95;
	ram[3724] = 8'h0c;	ram[3725] = 8'ha2;	ram[3726] = 8'h0e;	ram[3727] = 8'h47;
	ram[3728] = 8'h00;	ram[3729] = 8'h5f;	ram[3730] = 8'h0c;	ram[3731] = 8'hab;
	ram[3732] = 8'h0e;	ram[3733] = 8'h45;	ram[3734] = 8'h00;	ram[3735] = 8'h21;
	ram[3736] = 8'h0c;	ram[3737] = 8'h57;	ram[3738] = 8'h41;	ram[3739] = 8'h4e;
	ram[3740] = 8'h54;	ram[3741] = 8'h20;	ram[3742] = 8'h53;	ram[3743] = 8'h49;
	ram[3744] = 8'hce;	ram[3745] = 8'h00;	ram[3746] = 8'h57;	ram[3747] = 8'h41;
	ram[3748] = 8'h4e;	ram[3749] = 8'h54;	ram[3750] = 8'h20;	ram[3751] = 8'h52;
	ram[3752] = 8'h4e;	ram[3753] = 8'hc4;	ram[3754] = 8'h00;	ram[3755] = 8'h57;
	ram[3756] = 8'h41;	ram[3757] = 8'h4e;	ram[3758] = 8'h54;	ram[3759] = 8'h20;
	ram[3760] = 8'h53;	ram[3761] = 8'h51;	ram[3762] = 8'hd2;	ram[3763] = 8'h00;
	ram[3764] = 8'h54;	ram[3765] = 8'h45;	ram[3766] = 8'h52;	ram[3767] = 8'h4d;
	ram[3768] = 8'h49;	ram[3769] = 8'h4e;	ram[3770] = 8'h41;	ram[3771] = 8'h4c;
	ram[3772] = 8'h20;	ram[3773] = 8'h57;	ram[3774] = 8'h49;	ram[3775] = 8'h44;
	ram[3776] = 8'h54;	ram[3777] = 8'hc8;	ram[3778] = 8'h00;	ram[3779] = 8'h20;
	ram[3780] = 8'h42;	ram[3781] = 8'h59;	ram[3782] = 8'h54;	ram[3783] = 8'h45;
	ram[3784] = 8'h53;	ram[3785] = 8'h20;	ram[3786] = 8'h46;	ram[3787] = 8'h52;
	ram[3788] = 8'h45;	ram[3789] = 8'hc5;	ram[3790] = 8'h0d;	ram[3791] = 8'h0d;
	ram[3792] = 8'h42;	ram[3793] = 8'h41;	ram[3794] = 8'h53;	ram[3795] = 8'h49;
	ram[3796] = 8'h43;	ram[3797] = 8'h20;	ram[3798] = 8'h56;	ram[3799] = 8'h45;
	ram[3800] = 8'h52;	ram[3801] = 8'h53;	ram[3802] = 8'h49;	ram[3803] = 8'h4f;
	ram[3804] = 8'h4e;	ram[3805] = 8'h20;	ram[3806] = 8'h33;	ram[3807] = 8'h2e;
	ram[3808] = 8'hb2;	ram[3809] = 8'h0d;	ram[3810] = 8'h5b;	ram[3811] = 8'h34;
	ram[3812] = 8'h4b;	ram[3813] = 8'h20;	ram[3814] = 8'h56;	ram[3815] = 8'h45;
	ram[3816] = 8'h52;	ram[3817] = 8'h53;	ram[3818] = 8'h49;	ram[3819] = 8'h4f;
	ram[3820] = 8'h4e;	ram[3821] = 8'hdd;	ram[3822] = 8'h0d;	ram[3823] = 8'h00;
	ram[3824] = 8'h4d;	ram[3825] = 8'h45;	ram[3826] = 8'h4d;	ram[3827] = 8'h4f;
	ram[3828] = 8'h52;	ram[3829] = 8'h59;	ram[3830] = 8'h20;	ram[3831] = 8'h53;
	ram[3832] = 8'h49;	ram[3833] = 8'h5a;	ram[3834] = 8'hc5;	ram[3835] = 8'h00;
	ram[3836] = 8'h00;	ram[3837] = 8'h00;	ram[3838] = 8'h00;	ram[3839] = 8'h00;
	ram[3840] = 8'h00;	ram[3841] = 8'h00;	ram[3842] = 8'h00;	ram[3843] = 8'h00;
	ram[3844] = 8'h00;	ram[3845] = 8'h00;	ram[3846] = 8'h00;	ram[3847] = 8'h00;
	ram[3848] = 8'h00;	ram[3849] = 8'h00;	ram[3850] = 8'h00;	ram[3851] = 8'h00;
	ram[3852] = 8'h00;	ram[3853] = 8'h00;	ram[3854] = 8'h00;	ram[3855] = 8'h00;
	ram[3856] = 8'h00;	ram[3857] = 8'h00;	ram[3858] = 8'h00;	ram[3859] = 8'h00;
	ram[3860] = 8'h00;	ram[3861] = 8'h00;	ram[3862] = 8'h00;	ram[3863] = 8'h00;
	ram[3864] = 8'h00;	ram[3865] = 8'h00;	ram[3866] = 8'h00;	ram[3867] = 8'h00;
	ram[3868] = 8'h00;	ram[3869] = 8'h00;	ram[3870] = 8'h00;	ram[3871] = 8'h00;
	ram[3872] = 8'h00;	ram[3873] = 8'h00;	ram[3874] = 8'h00;	ram[3875] = 8'h00;
	ram[3876] = 8'h00;	ram[3877] = 8'h00;	ram[3878] = 8'h00;	ram[3879] = 8'h00;
	ram[3880] = 8'h00;	ram[3881] = 8'h00;	ram[3882] = 8'h00;	ram[3883] = 8'h00;
	ram[3884] = 8'h00;	ram[3885] = 8'h00;	ram[3886] = 8'h00;	ram[3887] = 8'h00;
	ram[3888] = 8'h00;	ram[3889] = 8'h00;	ram[3890] = 8'h00;	ram[3891] = 8'h00;
	ram[3892] = 8'h00;	ram[3893] = 8'h00;	ram[3894] = 8'h00;	ram[3895] = 8'h00;
	ram[3896] = 8'h00;	ram[3897] = 8'h00;	ram[3898] = 8'h00;	ram[3899] = 8'h00;
	ram[3900] = 8'h00;	ram[3901] = 8'h00;	ram[3902] = 8'h00;	ram[3903] = 8'h00;
	ram[3904] = 8'h00;	ram[3905] = 8'h00;	ram[3906] = 8'h00;	ram[3907] = 8'h00;
	ram[3908] = 8'h00;	ram[3909] = 8'h00;	ram[3910] = 8'h00;	ram[3911] = 8'h00;
	ram[3912] = 8'h00;	ram[3913] = 8'h00;	ram[3914] = 8'h00;	ram[3915] = 8'h00;
	ram[3916] = 8'h00;	ram[3917] = 8'h00;	ram[3918] = 8'h00;	ram[3919] = 8'h00;
	ram[3920] = 8'h00;	ram[3921] = 8'h00;	ram[3922] = 8'h00;	ram[3923] = 8'h00;
	ram[3924] = 8'h00;	ram[3925] = 8'h00;	ram[3926] = 8'h00;	ram[3927] = 8'h00;
	ram[3928] = 8'h00;	ram[3929] = 8'h00;	ram[3930] = 8'h00;	ram[3931] = 8'h00;
	ram[3932] = 8'h00;	ram[3933] = 8'h00;	ram[3934] = 8'h00;	ram[3935] = 8'h00;
	ram[3936] = 8'h00;	ram[3937] = 8'h00;	ram[3938] = 8'h00;	ram[3939] = 8'h00;
	ram[3940] = 8'h00;	ram[3941] = 8'h00;	ram[3942] = 8'h00;	ram[3943] = 8'h00;
	ram[3944] = 8'h00;	ram[3945] = 8'h00;	ram[3946] = 8'h00;	ram[3947] = 8'h00;
	ram[3948] = 8'h00;	ram[3949] = 8'h00;	ram[3950] = 8'h00;	ram[3951] = 8'h00;
	ram[3952] = 8'h00;	ram[3953] = 8'h00;	ram[3954] = 8'h00;	ram[3955] = 8'h00;
	ram[3956] = 8'h00;	ram[3957] = 8'h00;	ram[3958] = 8'h00;	ram[3959] = 8'h00;
	ram[3960] = 8'h00;	ram[3961] = 8'h00;	ram[3962] = 8'h00;	ram[3963] = 8'h00;
	ram[3964] = 8'h00;	ram[3965] = 8'h00;	ram[3966] = 8'h00;	ram[3967] = 8'h00;
	ram[3968] = 8'h00;	ram[3969] = 8'h00;	ram[3970] = 8'h00;	ram[3971] = 8'h00;
	ram[3972] = 8'h00;	ram[3973] = 8'h00;	ram[3974] = 8'h00;	ram[3975] = 8'h00;
	ram[3976] = 8'h00;	ram[3977] = 8'h00;	ram[3978] = 8'h00;	ram[3979] = 8'h00;
	ram[3980] = 8'h00;	ram[3981] = 8'h00;	ram[3982] = 8'h00;	ram[3983] = 8'h00;
	ram[3984] = 8'h00;	ram[3985] = 8'h00;	ram[3986] = 8'h00;	ram[3987] = 8'h00;
	ram[3988] = 8'h00;	ram[3989] = 8'h00;	ram[3990] = 8'h00;	ram[3991] = 8'h00;
	ram[3992] = 8'h00;	ram[3993] = 8'h00;	ram[3994] = 8'h00;	ram[3995] = 8'h00;
	ram[3996] = 8'h00;	ram[3997] = 8'h00;	ram[3998] = 8'h00;	ram[3999] = 8'h00;
	ram[4000] = 8'h00;	ram[4001] = 8'h00;	ram[4002] = 8'h00;	ram[4003] = 8'h00;
	ram[4004] = 8'h00;	ram[4005] = 8'h00;	ram[4006] = 8'h00;	ram[4007] = 8'h00;
	ram[4008] = 8'h00;	ram[4009] = 8'h00;	ram[4010] = 8'h00;	ram[4011] = 8'h00;
	ram[4012] = 8'h00;	ram[4013] = 8'h00;	ram[4014] = 8'h00;	ram[4015] = 8'h00;
	ram[4016] = 8'h00;	ram[4017] = 8'h00;	ram[4018] = 8'h00;	ram[4019] = 8'h00;
	ram[4020] = 8'h00;	ram[4021] = 8'h00;	ram[4022] = 8'h00;	ram[4023] = 8'h00;
	ram[4024] = 8'h00;	ram[4025] = 8'h00;	ram[4026] = 8'h00;	ram[4027] = 8'h00;
	ram[4028] = 8'h00;	ram[4029] = 8'h00;	ram[4030] = 8'h00;	ram[4031] = 8'h00;
	ram[4032] = 8'h00;	ram[4033] = 8'h00;	ram[4034] = 8'h00;	ram[4035] = 8'h00;
	ram[4036] = 8'h00;	ram[4037] = 8'h00;	ram[4038] = 8'h00;	ram[4039] = 8'h00;
	ram[4040] = 8'h00;	ram[4041] = 8'h00;	ram[4042] = 8'h00;	ram[4043] = 8'h00;
	ram[4044] = 8'h00;	ram[4045] = 8'h00;	ram[4046] = 8'h00;	ram[4047] = 8'h00;
	ram[4048] = 8'h00;	ram[4049] = 8'h00;	ram[4050] = 8'h00;	ram[4051] = 8'h00;
	ram[4052] = 8'h00;	ram[4053] = 8'h00;	ram[4054] = 8'h00;	ram[4055] = 8'h00;
	ram[4056] = 8'h00;	ram[4057] = 8'h00;	ram[4058] = 8'h00;	ram[4059] = 8'h00;
	ram[4060] = 8'h00;	ram[4061] = 8'h00;	ram[4062] = 8'h00;	ram[4063] = 8'h00;
	ram[4064] = 8'h00;	ram[4065] = 8'h00;	ram[4066] = 8'h00;	ram[4067] = 8'h00;
	ram[4068] = 8'h00;	ram[4069] = 8'h00;	ram[4070] = 8'h00;	ram[4071] = 8'h00;
	ram[4072] = 8'h00;	ram[4073] = 8'h00;	ram[4074] = 8'h00;	ram[4075] = 8'h00;
	ram[4076] = 8'h00;	ram[4077] = 8'h00;	ram[4078] = 8'h00;	ram[4079] = 8'h00;
	ram[4080] = 8'h00;	ram[4081] = 8'h00;	ram[4082] = 8'h00;	ram[4083] = 8'h00;
	ram[4084] = 8'h00;	ram[4085] = 8'h00;	ram[4086] = 8'h00;	ram[4087] = 8'h00;
	ram[4088] = 8'h00;	ram[4089] = 8'h00;	ram[4090] = 8'h00;	ram[4091] = 8'h00;
	ram[4092] = 8'h00;	ram[4093] = 8'h00;	ram[4094] = 8'h00;	ram[4095] = 8'h00;
	ram[4096] = 8'h00;	ram[4097] = 8'h00;	ram[4098] = 8'h00;	ram[4099] = 8'h00;
	ram[4100] = 8'h00;	ram[4101] = 8'h00;	ram[4102] = 8'h00;	ram[4103] = 8'h00;
	ram[4104] = 8'h00;	ram[4105] = 8'h00;	ram[4106] = 8'h00;	ram[4107] = 8'h00;
	ram[4108] = 8'h00;	ram[4109] = 8'h00;	ram[4110] = 8'h00;	ram[4111] = 8'h00;
	ram[4112] = 8'h00;	ram[4113] = 8'h00;	ram[4114] = 8'h00;	ram[4115] = 8'h00;
	ram[4116] = 8'h00;	ram[4117] = 8'h00;	ram[4118] = 8'h00;	ram[4119] = 8'h00;
	ram[4120] = 8'h00;	ram[4121] = 8'h00;	ram[4122] = 8'h00;	ram[4123] = 8'h00;
	ram[4124] = 8'h00;	ram[4125] = 8'h00;	ram[4126] = 8'h00;	ram[4127] = 8'h00;
	ram[4128] = 8'h00;	ram[4129] = 8'h00;	ram[4130] = 8'h00;	ram[4131] = 8'h00;
	ram[4132] = 8'h00;	ram[4133] = 8'h00;	ram[4134] = 8'h00;	ram[4135] = 8'h00;
	ram[4136] = 8'h00;	ram[4137] = 8'h00;	ram[4138] = 8'h00;	ram[4139] = 8'h00;
	ram[4140] = 8'h00;	ram[4141] = 8'h00;	ram[4142] = 8'h00;	ram[4143] = 8'h00;
	ram[4144] = 8'h00;	ram[4145] = 8'h00;	ram[4146] = 8'h00;	ram[4147] = 8'h00;
	ram[4148] = 8'h00;	ram[4149] = 8'h00;	ram[4150] = 8'h00;	ram[4151] = 8'h00;
	ram[4152] = 8'h00;	ram[4153] = 8'h00;	ram[4154] = 8'h00;	ram[4155] = 8'h00;
	ram[4156] = 8'h00;	ram[4157] = 8'h00;	ram[4158] = 8'h00;	ram[4159] = 8'h00;
	ram[4160] = 8'h00;	ram[4161] = 8'h00;	ram[4162] = 8'h00;	ram[4163] = 8'h00;
	ram[4164] = 8'h00;	ram[4165] = 8'h00;	ram[4166] = 8'h00;	ram[4167] = 8'h00;
	ram[4168] = 8'h00;	ram[4169] = 8'h00;	ram[4170] = 8'h00;	ram[4171] = 8'h00;
	ram[4172] = 8'h00;	ram[4173] = 8'h00;	ram[4174] = 8'h00;	ram[4175] = 8'h00;
	ram[4176] = 8'h00;	ram[4177] = 8'h00;	ram[4178] = 8'h00;	ram[4179] = 8'h00;
	ram[4180] = 8'h00;	ram[4181] = 8'h00;	ram[4182] = 8'h00;	ram[4183] = 8'h00;
	ram[4184] = 8'h00;	ram[4185] = 8'h00;	ram[4186] = 8'h00;	ram[4187] = 8'h00;
	ram[4188] = 8'h00;	ram[4189] = 8'h00;	ram[4190] = 8'h00;	ram[4191] = 8'h00;
	ram[4192] = 8'h00;	ram[4193] = 8'h00;	ram[4194] = 8'h00;	ram[4195] = 8'h00;
	ram[4196] = 8'h00;	ram[4197] = 8'h00;	ram[4198] = 8'h00;	ram[4199] = 8'h00;
	ram[4200] = 8'h00;	ram[4201] = 8'h00;	ram[4202] = 8'h00;	ram[4203] = 8'h00;
	ram[4204] = 8'h00;	ram[4205] = 8'h00;	ram[4206] = 8'h00;	ram[4207] = 8'h00;
	ram[4208] = 8'h00;	ram[4209] = 8'h00;	ram[4210] = 8'h00;	ram[4211] = 8'h00;
	ram[4212] = 8'h00;	ram[4213] = 8'h00;	ram[4214] = 8'h00;	ram[4215] = 8'h00;
	ram[4216] = 8'h00;	ram[4217] = 8'h00;	ram[4218] = 8'h00;	ram[4219] = 8'h00;
	ram[4220] = 8'h00;	ram[4221] = 8'h00;	ram[4222] = 8'h00;	ram[4223] = 8'h00;
	ram[4224] = 8'h00;	ram[4225] = 8'h00;	ram[4226] = 8'h00;	ram[4227] = 8'h00;
	ram[4228] = 8'h00;	ram[4229] = 8'h00;	ram[4230] = 8'h00;	ram[4231] = 8'h00;
	ram[4232] = 8'h00;	ram[4233] = 8'h00;	ram[4234] = 8'h00;	ram[4235] = 8'h00;
	ram[4236] = 8'h00;	ram[4237] = 8'h00;	ram[4238] = 8'h00;	ram[4239] = 8'h00;
	ram[4240] = 8'h00;	ram[4241] = 8'h00;	ram[4242] = 8'h00;	ram[4243] = 8'h00;
	ram[4244] = 8'h00;	ram[4245] = 8'h00;	ram[4246] = 8'h00;	ram[4247] = 8'h00;
	ram[4248] = 8'h00;	ram[4249] = 8'h00;	ram[4250] = 8'h00;	ram[4251] = 8'h00;
	ram[4252] = 8'h00;	ram[4253] = 8'h00;	ram[4254] = 8'h00;	ram[4255] = 8'h00;
	ram[4256] = 8'h00;	ram[4257] = 8'h00;	ram[4258] = 8'h00;	ram[4259] = 8'h00;
	ram[4260] = 8'h00;	ram[4261] = 8'h00;	ram[4262] = 8'h00;	ram[4263] = 8'h00;
	ram[4264] = 8'h00;	ram[4265] = 8'h00;	ram[4266] = 8'h00;	ram[4267] = 8'h00;
	ram[4268] = 8'h00;	ram[4269] = 8'h00;	ram[4270] = 8'h00;	ram[4271] = 8'h00;
	ram[4272] = 8'h00;	ram[4273] = 8'h00;	ram[4274] = 8'h00;	ram[4275] = 8'h00;
	ram[4276] = 8'h00;	ram[4277] = 8'h00;	ram[4278] = 8'h00;	ram[4279] = 8'h00;
	ram[4280] = 8'h00;	ram[4281] = 8'h00;	ram[4282] = 8'h00;	ram[4283] = 8'h00;
	ram[4284] = 8'h00;	ram[4285] = 8'h00;	ram[4286] = 8'h00;	ram[4287] = 8'h00;
	ram[4288] = 8'h00;	ram[4289] = 8'h00;	ram[4290] = 8'h00;	ram[4291] = 8'h00;
	ram[4292] = 8'h00;	ram[4293] = 8'h00;	ram[4294] = 8'h00;	ram[4295] = 8'h00;
	ram[4296] = 8'h00;	ram[4297] = 8'h00;	ram[4298] = 8'h00;	ram[4299] = 8'h00;
	ram[4300] = 8'h00;	ram[4301] = 8'h00;	ram[4302] = 8'h00;	ram[4303] = 8'h00;
	ram[4304] = 8'h00;	ram[4305] = 8'h00;	ram[4306] = 8'h00;	ram[4307] = 8'h00;
	ram[4308] = 8'h00;	ram[4309] = 8'h00;	ram[4310] = 8'h00;	ram[4311] = 8'h00;
	ram[4312] = 8'h00;	ram[4313] = 8'h00;	ram[4314] = 8'h00;	ram[4315] = 8'h00;
	ram[4316] = 8'h00;	ram[4317] = 8'h00;	ram[4318] = 8'h00;	ram[4319] = 8'h00;
	ram[4320] = 8'h00;	ram[4321] = 8'h00;	ram[4322] = 8'h00;	ram[4323] = 8'h00;
	ram[4324] = 8'h00;	ram[4325] = 8'h00;	ram[4326] = 8'h00;	ram[4327] = 8'h00;
	ram[4328] = 8'h00;	ram[4329] = 8'h00;	ram[4330] = 8'h00;	ram[4331] = 8'h00;
	ram[4332] = 8'h00;	ram[4333] = 8'h00;	ram[4334] = 8'h00;	ram[4335] = 8'h00;
	ram[4336] = 8'h00;	ram[4337] = 8'h00;	ram[4338] = 8'h00;	ram[4339] = 8'h00;
	ram[4340] = 8'h00;	ram[4341] = 8'h00;	ram[4342] = 8'h00;	ram[4343] = 8'h00;
	ram[4344] = 8'h00;	ram[4345] = 8'h00;	ram[4346] = 8'h00;	ram[4347] = 8'h00;
	ram[4348] = 8'h00;	ram[4349] = 8'h00;	ram[4350] = 8'h00;	ram[4351] = 8'h00;
	ram[4352] = 8'h00;	ram[4353] = 8'h00;	ram[4354] = 8'h00;	ram[4355] = 8'h00;
	ram[4356] = 8'h00;	ram[4357] = 8'h00;	ram[4358] = 8'h00;	ram[4359] = 8'h00;
	ram[4360] = 8'h00;	ram[4361] = 8'h00;	ram[4362] = 8'h00;	ram[4363] = 8'h00;
	ram[4364] = 8'h00;	ram[4365] = 8'h00;	ram[4366] = 8'h00;	ram[4367] = 8'h00;
	ram[4368] = 8'h00;	ram[4369] = 8'h00;	ram[4370] = 8'h00;	ram[4371] = 8'h00;
	ram[4372] = 8'h00;	ram[4373] = 8'h00;	ram[4374] = 8'h00;	ram[4375] = 8'h00;
	ram[4376] = 8'h00;	ram[4377] = 8'h00;	ram[4378] = 8'h00;	ram[4379] = 8'h00;
	ram[4380] = 8'h00;	ram[4381] = 8'h00;	ram[4382] = 8'h00;	ram[4383] = 8'h00;
	ram[4384] = 8'h00;	ram[4385] = 8'h00;	ram[4386] = 8'h00;	ram[4387] = 8'h00;
	ram[4388] = 8'h00;	ram[4389] = 8'h00;	ram[4390] = 8'h00;	ram[4391] = 8'h00;
	ram[4392] = 8'h00;	ram[4393] = 8'h00;	ram[4394] = 8'h00;	ram[4395] = 8'h00;
	ram[4396] = 8'h00;	ram[4397] = 8'h00;	ram[4398] = 8'h00;	ram[4399] = 8'h00;
	ram[4400] = 8'h00;	ram[4401] = 8'h00;	ram[4402] = 8'h00;	ram[4403] = 8'h00;
	ram[4404] = 8'h00;	ram[4405] = 8'h00;	ram[4406] = 8'h00;	ram[4407] = 8'h00;
	ram[4408] = 8'h00;	ram[4409] = 8'h00;	ram[4410] = 8'h00;	ram[4411] = 8'h00;
	ram[4412] = 8'h00;	ram[4413] = 8'h00;	ram[4414] = 8'h00;	ram[4415] = 8'h00;
	ram[4416] = 8'h00;	ram[4417] = 8'h00;	ram[4418] = 8'h00;	ram[4419] = 8'h00;
	ram[4420] = 8'h00;	ram[4421] = 8'h00;	ram[4422] = 8'h00;	ram[4423] = 8'h00;
	ram[4424] = 8'h00;	ram[4425] = 8'h00;	ram[4426] = 8'h00;	ram[4427] = 8'h00;
	ram[4428] = 8'h00;	ram[4429] = 8'h00;	ram[4430] = 8'h00;	ram[4431] = 8'h00;
	ram[4432] = 8'h00;	ram[4433] = 8'h00;	ram[4434] = 8'h00;	ram[4435] = 8'h00;
	ram[4436] = 8'h00;	ram[4437] = 8'h00;	ram[4438] = 8'h00;	ram[4439] = 8'h00;
	ram[4440] = 8'h00;	ram[4441] = 8'h00;	ram[4442] = 8'h00;	ram[4443] = 8'h00;
	ram[4444] = 8'h00;	ram[4445] = 8'h00;	ram[4446] = 8'h00;	ram[4447] = 8'h00;
	ram[4448] = 8'h00;	ram[4449] = 8'h00;	ram[4450] = 8'h00;	ram[4451] = 8'h00;
	ram[4452] = 8'h00;	ram[4453] = 8'h00;	ram[4454] = 8'h00;	ram[4455] = 8'h00;
	ram[4456] = 8'h00;	ram[4457] = 8'h00;	ram[4458] = 8'h00;	ram[4459] = 8'h00;
	ram[4460] = 8'h00;	ram[4461] = 8'h00;	ram[4462] = 8'h00;	ram[4463] = 8'h00;
	ram[4464] = 8'h00;	ram[4465] = 8'h00;	ram[4466] = 8'h00;	ram[4467] = 8'h00;
	ram[4468] = 8'h00;	ram[4469] = 8'h00;	ram[4470] = 8'h00;	ram[4471] = 8'h00;
	ram[4472] = 8'h00;	ram[4473] = 8'h00;	ram[4474] = 8'h00;	ram[4475] = 8'h00;
	ram[4476] = 8'h00;	ram[4477] = 8'h00;	ram[4478] = 8'h00;	ram[4479] = 8'h00;
	ram[4480] = 8'h00;	ram[4481] = 8'h00;	ram[4482] = 8'h00;	ram[4483] = 8'h00;
	ram[4484] = 8'h00;	ram[4485] = 8'h00;	ram[4486] = 8'h00;	ram[4487] = 8'h00;
	ram[4488] = 8'h00;	ram[4489] = 8'h00;	ram[4490] = 8'h00;	ram[4491] = 8'h00;
	ram[4492] = 8'h00;	ram[4493] = 8'h00;	ram[4494] = 8'h00;	ram[4495] = 8'h00;
	ram[4496] = 8'h00;	ram[4497] = 8'h00;	ram[4498] = 8'h00;	ram[4499] = 8'h00;
	ram[4500] = 8'h00;	ram[4501] = 8'h00;	ram[4502] = 8'h00;	ram[4503] = 8'h00;
	ram[4504] = 8'h00;	ram[4505] = 8'h00;	ram[4506] = 8'h00;	ram[4507] = 8'h00;
	ram[4508] = 8'h00;	ram[4509] = 8'h00;	ram[4510] = 8'h00;	ram[4511] = 8'h00;
	ram[4512] = 8'h00;	ram[4513] = 8'h00;	ram[4514] = 8'h00;	ram[4515] = 8'h00;
	ram[4516] = 8'h00;	ram[4517] = 8'h00;	ram[4518] = 8'h00;	ram[4519] = 8'h00;
	ram[4520] = 8'h00;	ram[4521] = 8'h00;	ram[4522] = 8'h00;	ram[4523] = 8'h00;
	ram[4524] = 8'h00;	ram[4525] = 8'h00;	ram[4526] = 8'h00;	ram[4527] = 8'h00;
	ram[4528] = 8'h00;	ram[4529] = 8'h00;	ram[4530] = 8'h00;	ram[4531] = 8'h00;
	ram[4532] = 8'h00;	ram[4533] = 8'h00;	ram[4534] = 8'h00;	ram[4535] = 8'h00;
	ram[4536] = 8'h00;	ram[4537] = 8'h00;	ram[4538] = 8'h00;	ram[4539] = 8'h00;
	ram[4540] = 8'h00;	ram[4541] = 8'h00;	ram[4542] = 8'h00;	ram[4543] = 8'h00;
	ram[4544] = 8'h00;	ram[4545] = 8'h00;	ram[4546] = 8'h00;	ram[4547] = 8'h00;
	ram[4548] = 8'h00;	ram[4549] = 8'h00;	ram[4550] = 8'h00;	ram[4551] = 8'h00;
	ram[4552] = 8'h00;	ram[4553] = 8'h00;	ram[4554] = 8'h00;	ram[4555] = 8'h00;
	ram[4556] = 8'h00;	ram[4557] = 8'h00;	ram[4558] = 8'h00;	ram[4559] = 8'h00;
	ram[4560] = 8'h00;	ram[4561] = 8'h00;	ram[4562] = 8'h00;	ram[4563] = 8'h00;
	ram[4564] = 8'h00;	ram[4565] = 8'h00;	ram[4566] = 8'h00;	ram[4567] = 8'h00;
	ram[4568] = 8'h00;	ram[4569] = 8'h00;	ram[4570] = 8'h00;	ram[4571] = 8'h00;
	ram[4572] = 8'h00;	ram[4573] = 8'h00;	ram[4574] = 8'h00;	ram[4575] = 8'h00;
	ram[4576] = 8'h00;	ram[4577] = 8'h00;	ram[4578] = 8'h00;	ram[4579] = 8'h00;
	ram[4580] = 8'h00;	ram[4581] = 8'h00;	ram[4582] = 8'h00;	ram[4583] = 8'h00;
	ram[4584] = 8'h00;	ram[4585] = 8'h00;	ram[4586] = 8'h00;	ram[4587] = 8'h00;
	ram[4588] = 8'h00;	ram[4589] = 8'h00;	ram[4590] = 8'h00;	ram[4591] = 8'h00;
	ram[4592] = 8'h00;	ram[4593] = 8'h00;	ram[4594] = 8'h00;	ram[4595] = 8'h00;
	ram[4596] = 8'h00;	ram[4597] = 8'h00;	ram[4598] = 8'h00;	ram[4599] = 8'h00;
	ram[4600] = 8'h00;	ram[4601] = 8'h00;	ram[4602] = 8'h00;	ram[4603] = 8'h00;
	ram[4604] = 8'h00;	ram[4605] = 8'h00;	ram[4606] = 8'h00;	ram[4607] = 8'h00;
	ram[4608] = 8'h00;	ram[4609] = 8'h00;	ram[4610] = 8'h00;	ram[4611] = 8'h00;
	ram[4612] = 8'h00;	ram[4613] = 8'h00;	ram[4614] = 8'h00;	ram[4615] = 8'h00;
	ram[4616] = 8'h00;	ram[4617] = 8'h00;	ram[4618] = 8'h00;	ram[4619] = 8'h00;
	ram[4620] = 8'h00;	ram[4621] = 8'h00;	ram[4622] = 8'h00;	ram[4623] = 8'h00;
	ram[4624] = 8'h00;	ram[4625] = 8'h00;	ram[4626] = 8'h00;	ram[4627] = 8'h00;
	ram[4628] = 8'h00;	ram[4629] = 8'h00;	ram[4630] = 8'h00;	ram[4631] = 8'h00;
	ram[4632] = 8'h00;	ram[4633] = 8'h00;	ram[4634] = 8'h00;	ram[4635] = 8'h00;
	ram[4636] = 8'h00;	ram[4637] = 8'h00;	ram[4638] = 8'h00;	ram[4639] = 8'h00;
	ram[4640] = 8'h00;	ram[4641] = 8'h00;	ram[4642] = 8'h00;	ram[4643] = 8'h00;
	ram[4644] = 8'h00;	ram[4645] = 8'h00;	ram[4646] = 8'h00;	ram[4647] = 8'h00;
	ram[4648] = 8'h00;	ram[4649] = 8'h00;	ram[4650] = 8'h00;	ram[4651] = 8'h00;
	ram[4652] = 8'h00;	ram[4653] = 8'h00;	ram[4654] = 8'h00;	ram[4655] = 8'h00;
	ram[4656] = 8'h00;	ram[4657] = 8'h00;	ram[4658] = 8'h00;	ram[4659] = 8'h00;
	ram[4660] = 8'h00;	ram[4661] = 8'h00;	ram[4662] = 8'h00;	ram[4663] = 8'h00;
	ram[4664] = 8'h00;	ram[4665] = 8'h00;	ram[4666] = 8'h00;	ram[4667] = 8'h00;
	ram[4668] = 8'h00;	ram[4669] = 8'h00;	ram[4670] = 8'h00;	ram[4671] = 8'h00;
	ram[4672] = 8'h00;	ram[4673] = 8'h00;	ram[4674] = 8'h00;	ram[4675] = 8'h00;
	ram[4676] = 8'h00;	ram[4677] = 8'h00;	ram[4678] = 8'h00;	ram[4679] = 8'h00;
	ram[4680] = 8'h00;	ram[4681] = 8'h00;	ram[4682] = 8'h00;	ram[4683] = 8'h00;
	ram[4684] = 8'h00;	ram[4685] = 8'h00;	ram[4686] = 8'h00;	ram[4687] = 8'h00;
	ram[4688] = 8'h00;	ram[4689] = 8'h00;	ram[4690] = 8'h00;	ram[4691] = 8'h00;
	ram[4692] = 8'h00;	ram[4693] = 8'h00;	ram[4694] = 8'h00;	ram[4695] = 8'h00;
	ram[4696] = 8'h00;	ram[4697] = 8'h00;	ram[4698] = 8'h00;	ram[4699] = 8'h00;
	ram[4700] = 8'h00;	ram[4701] = 8'h00;	ram[4702] = 8'h00;	ram[4703] = 8'h00;
	ram[4704] = 8'h00;	ram[4705] = 8'h00;	ram[4706] = 8'h00;	ram[4707] = 8'h00;
	ram[4708] = 8'h00;	ram[4709] = 8'h00;	ram[4710] = 8'h00;	ram[4711] = 8'h00;
	ram[4712] = 8'h00;	ram[4713] = 8'h00;	ram[4714] = 8'h00;	ram[4715] = 8'h00;
	ram[4716] = 8'h00;	ram[4717] = 8'h00;	ram[4718] = 8'h00;	ram[4719] = 8'h00;
	ram[4720] = 8'h00;	ram[4721] = 8'h00;	ram[4722] = 8'h00;	ram[4723] = 8'h00;
	ram[4724] = 8'h00;	ram[4725] = 8'h00;	ram[4726] = 8'h00;	ram[4727] = 8'h00;
	ram[4728] = 8'h00;	ram[4729] = 8'h00;	ram[4730] = 8'h00;	ram[4731] = 8'h00;
	ram[4732] = 8'h00;	ram[4733] = 8'h00;	ram[4734] = 8'h00;	ram[4735] = 8'h00;
	ram[4736] = 8'h00;	ram[4737] = 8'h00;	ram[4738] = 8'h00;	ram[4739] = 8'h00;
	ram[4740] = 8'h00;	ram[4741] = 8'h00;	ram[4742] = 8'h00;	ram[4743] = 8'h00;
	ram[4744] = 8'h00;	ram[4745] = 8'h00;	ram[4746] = 8'h00;	ram[4747] = 8'h00;
	ram[4748] = 8'h00;	ram[4749] = 8'h00;	ram[4750] = 8'h00;	ram[4751] = 8'h00;
	ram[4752] = 8'h00;	ram[4753] = 8'h00;	ram[4754] = 8'h00;	ram[4755] = 8'h00;
	ram[4756] = 8'h00;	ram[4757] = 8'h00;	ram[4758] = 8'h00;	ram[4759] = 8'h00;
	ram[4760] = 8'h00;	ram[4761] = 8'h00;	ram[4762] = 8'h00;	ram[4763] = 8'h00;
	ram[4764] = 8'h00;	ram[4765] = 8'h00;	ram[4766] = 8'h00;	ram[4767] = 8'h00;
	ram[4768] = 8'h00;	ram[4769] = 8'h00;	ram[4770] = 8'h00;	ram[4771] = 8'h00;
	ram[4772] = 8'h00;	ram[4773] = 8'h00;	ram[4774] = 8'h00;	ram[4775] = 8'h00;
	ram[4776] = 8'h00;	ram[4777] = 8'h00;	ram[4778] = 8'h00;	ram[4779] = 8'h00;
	ram[4780] = 8'h00;	ram[4781] = 8'h00;	ram[4782] = 8'h00;	ram[4783] = 8'h00;
	ram[4784] = 8'h00;	ram[4785] = 8'h00;	ram[4786] = 8'h00;	ram[4787] = 8'h00;
	ram[4788] = 8'h00;	ram[4789] = 8'h00;	ram[4790] = 8'h00;	ram[4791] = 8'h00;
	ram[4792] = 8'h00;	ram[4793] = 8'h00;	ram[4794] = 8'h00;	ram[4795] = 8'h00;
	ram[4796] = 8'h00;	ram[4797] = 8'h00;	ram[4798] = 8'h00;	ram[4799] = 8'h00;
	ram[4800] = 8'h00;	ram[4801] = 8'h00;	ram[4802] = 8'h00;	ram[4803] = 8'h00;
	ram[4804] = 8'h00;	ram[4805] = 8'h00;	ram[4806] = 8'h00;	ram[4807] = 8'h00;
	ram[4808] = 8'h00;	ram[4809] = 8'h00;	ram[4810] = 8'h00;	ram[4811] = 8'h00;
	ram[4812] = 8'h00;	ram[4813] = 8'h00;	ram[4814] = 8'h00;	ram[4815] = 8'h00;
	ram[4816] = 8'h00;	ram[4817] = 8'h00;	ram[4818] = 8'h00;	ram[4819] = 8'h00;
	ram[4820] = 8'h00;	ram[4821] = 8'h00;	ram[4822] = 8'h00;	ram[4823] = 8'h00;
	ram[4824] = 8'h00;	ram[4825] = 8'h00;	ram[4826] = 8'h00;	ram[4827] = 8'h00;
	ram[4828] = 8'h00;	ram[4829] = 8'h00;	ram[4830] = 8'h00;	ram[4831] = 8'h00;
	ram[4832] = 8'h00;	ram[4833] = 8'h00;	ram[4834] = 8'h00;	ram[4835] = 8'h00;
	ram[4836] = 8'h00;	ram[4837] = 8'h00;	ram[4838] = 8'h00;	ram[4839] = 8'h00;
	ram[4840] = 8'h00;	ram[4841] = 8'h00;	ram[4842] = 8'h00;	ram[4843] = 8'h00;
	ram[4844] = 8'h00;	ram[4845] = 8'h00;	ram[4846] = 8'h00;	ram[4847] = 8'h00;
	ram[4848] = 8'h00;	ram[4849] = 8'h00;	ram[4850] = 8'h00;	ram[4851] = 8'h00;
	ram[4852] = 8'h00;	ram[4853] = 8'h00;	ram[4854] = 8'h00;	ram[4855] = 8'h00;
	ram[4856] = 8'h00;	ram[4857] = 8'h00;	ram[4858] = 8'h00;	ram[4859] = 8'h00;
	ram[4860] = 8'h00;	ram[4861] = 8'h00;	ram[4862] = 8'h00;	ram[4863] = 8'h00;
	ram[4864] = 8'h00;	ram[4865] = 8'h00;	ram[4866] = 8'h00;	ram[4867] = 8'h00;
	ram[4868] = 8'h00;	ram[4869] = 8'h00;	ram[4870] = 8'h00;	ram[4871] = 8'h00;
	ram[4872] = 8'h00;	ram[4873] = 8'h00;	ram[4874] = 8'h00;	ram[4875] = 8'h00;
	ram[4876] = 8'h00;	ram[4877] = 8'h00;	ram[4878] = 8'h00;	ram[4879] = 8'h00;
	ram[4880] = 8'h00;	ram[4881] = 8'h00;	ram[4882] = 8'h00;	ram[4883] = 8'h00;
	ram[4884] = 8'h00;	ram[4885] = 8'h00;	ram[4886] = 8'h00;	ram[4887] = 8'h00;
	ram[4888] = 8'h00;	ram[4889] = 8'h00;	ram[4890] = 8'h00;	ram[4891] = 8'h00;
	ram[4892] = 8'h00;	ram[4893] = 8'h00;	ram[4894] = 8'h00;	ram[4895] = 8'h00;
	ram[4896] = 8'h00;	ram[4897] = 8'h00;	ram[4898] = 8'h00;	ram[4899] = 8'h00;
	ram[4900] = 8'h00;	ram[4901] = 8'h00;	ram[4902] = 8'h00;	ram[4903] = 8'h00;
	ram[4904] = 8'h00;	ram[4905] = 8'h00;	ram[4906] = 8'h00;	ram[4907] = 8'h00;
	ram[4908] = 8'h00;	ram[4909] = 8'h00;	ram[4910] = 8'h00;	ram[4911] = 8'h00;
	ram[4912] = 8'h00;	ram[4913] = 8'h00;	ram[4914] = 8'h00;	ram[4915] = 8'h00;
	ram[4916] = 8'h00;	ram[4917] = 8'h00;	ram[4918] = 8'h00;	ram[4919] = 8'h00;
	ram[4920] = 8'h00;	ram[4921] = 8'h00;	ram[4922] = 8'h00;	ram[4923] = 8'h00;
	ram[4924] = 8'h00;	ram[4925] = 8'h00;	ram[4926] = 8'h00;	ram[4927] = 8'h00;
	ram[4928] = 8'h00;	ram[4929] = 8'h00;	ram[4930] = 8'h00;	ram[4931] = 8'h00;
	ram[4932] = 8'h00;	ram[4933] = 8'h00;	ram[4934] = 8'h00;	ram[4935] = 8'h00;
	ram[4936] = 8'h00;	ram[4937] = 8'h00;	ram[4938] = 8'h00;	ram[4939] = 8'h00;
	ram[4940] = 8'h00;	ram[4941] = 8'h00;	ram[4942] = 8'h00;	ram[4943] = 8'h00;
	ram[4944] = 8'h00;	ram[4945] = 8'h00;	ram[4946] = 8'h00;	ram[4947] = 8'h00;
	ram[4948] = 8'h00;	ram[4949] = 8'h00;	ram[4950] = 8'h00;	ram[4951] = 8'h00;
	ram[4952] = 8'h00;	ram[4953] = 8'h00;	ram[4954] = 8'h00;	ram[4955] = 8'h00;
	ram[4956] = 8'h00;	ram[4957] = 8'h00;	ram[4958] = 8'h00;	ram[4959] = 8'h00;
	ram[4960] = 8'h00;	ram[4961] = 8'h00;	ram[4962] = 8'h00;	ram[4963] = 8'h00;
	ram[4964] = 8'h00;	ram[4965] = 8'h00;	ram[4966] = 8'h00;	ram[4967] = 8'h00;
	ram[4968] = 8'h00;	ram[4969] = 8'h00;	ram[4970] = 8'h00;	ram[4971] = 8'h00;
	ram[4972] = 8'h00;	ram[4973] = 8'h00;	ram[4974] = 8'h00;	ram[4975] = 8'h00;
	ram[4976] = 8'h00;	ram[4977] = 8'h00;	ram[4978] = 8'h00;	ram[4979] = 8'h00;
	ram[4980] = 8'h00;	ram[4981] = 8'h00;	ram[4982] = 8'h00;	ram[4983] = 8'h00;
	ram[4984] = 8'h00;	ram[4985] = 8'h00;	ram[4986] = 8'h00;	ram[4987] = 8'h00;
	ram[4988] = 8'h00;	ram[4989] = 8'h00;	ram[4990] = 8'h00;	ram[4991] = 8'h00;
	ram[4992] = 8'h00;	ram[4993] = 8'h00;	ram[4994] = 8'h00;	ram[4995] = 8'h00;
	ram[4996] = 8'h00;	ram[4997] = 8'h00;	ram[4998] = 8'h00;	ram[4999] = 8'h00;
	ram[5000] = 8'h00;	ram[5001] = 8'h00;	ram[5002] = 8'h00;	ram[5003] = 8'h00;
	ram[5004] = 8'h00;	ram[5005] = 8'h00;	ram[5006] = 8'h00;	ram[5007] = 8'h00;
	ram[5008] = 8'h00;	ram[5009] = 8'h00;	ram[5010] = 8'h00;	ram[5011] = 8'h00;
	ram[5012] = 8'h00;	ram[5013] = 8'h00;	ram[5014] = 8'h00;	ram[5015] = 8'h00;
	ram[5016] = 8'h00;	ram[5017] = 8'h00;	ram[5018] = 8'h00;	ram[5019] = 8'h00;
	ram[5020] = 8'h00;	ram[5021] = 8'h00;	ram[5022] = 8'h00;	ram[5023] = 8'h00;
	ram[5024] = 8'h00;	ram[5025] = 8'h00;	ram[5026] = 8'h00;	ram[5027] = 8'h00;
	ram[5028] = 8'h00;	ram[5029] = 8'h00;	ram[5030] = 8'h00;	ram[5031] = 8'h00;
	ram[5032] = 8'h00;	ram[5033] = 8'h00;	ram[5034] = 8'h00;	ram[5035] = 8'h00;
	ram[5036] = 8'h00;	ram[5037] = 8'h00;	ram[5038] = 8'h00;	ram[5039] = 8'h00;
	ram[5040] = 8'h00;	ram[5041] = 8'h00;	ram[5042] = 8'h00;	ram[5043] = 8'h00;
	ram[5044] = 8'h00;	ram[5045] = 8'h00;	ram[5046] = 8'h00;	ram[5047] = 8'h00;
	ram[5048] = 8'h00;	ram[5049] = 8'h00;	ram[5050] = 8'h00;	ram[5051] = 8'h00;
	ram[5052] = 8'h00;	ram[5053] = 8'h00;	ram[5054] = 8'h00;	ram[5055] = 8'h00;
	ram[5056] = 8'h00;	ram[5057] = 8'h00;	ram[5058] = 8'h00;	ram[5059] = 8'h00;
	ram[5060] = 8'h00;	ram[5061] = 8'h00;	ram[5062] = 8'h00;	ram[5063] = 8'h00;
	ram[5064] = 8'h00;	ram[5065] = 8'h00;	ram[5066] = 8'h00;	ram[5067] = 8'h00;
	ram[5068] = 8'h00;	ram[5069] = 8'h00;	ram[5070] = 8'h00;	ram[5071] = 8'h00;
	ram[5072] = 8'h00;	ram[5073] = 8'h00;	ram[5074] = 8'h00;	ram[5075] = 8'h00;
	ram[5076] = 8'h00;	ram[5077] = 8'h00;	ram[5078] = 8'h00;	ram[5079] = 8'h00;
	ram[5080] = 8'h00;	ram[5081] = 8'h00;	ram[5082] = 8'h00;	ram[5083] = 8'h00;
	ram[5084] = 8'h00;	ram[5085] = 8'h00;	ram[5086] = 8'h00;	ram[5087] = 8'h00;
	ram[5088] = 8'h00;	ram[5089] = 8'h00;	ram[5090] = 8'h00;	ram[5091] = 8'h00;
	ram[5092] = 8'h00;	ram[5093] = 8'h00;	ram[5094] = 8'h00;	ram[5095] = 8'h00;
	ram[5096] = 8'h00;	ram[5097] = 8'h00;	ram[5098] = 8'h00;	ram[5099] = 8'h00;
	ram[5100] = 8'h00;	ram[5101] = 8'h00;	ram[5102] = 8'h00;	ram[5103] = 8'h00;
	ram[5104] = 8'h00;	ram[5105] = 8'h00;	ram[5106] = 8'h00;	ram[5107] = 8'h00;
	ram[5108] = 8'h00;	ram[5109] = 8'h00;	ram[5110] = 8'h00;	ram[5111] = 8'h00;
	ram[5112] = 8'h00;	ram[5113] = 8'h00;	ram[5114] = 8'h00;	ram[5115] = 8'h00;
	ram[5116] = 8'h00;	ram[5117] = 8'h00;	ram[5118] = 8'h00;	ram[5119] = 8'h00;
	ram[5120] = 8'h00;	ram[5121] = 8'h00;	ram[5122] = 8'h00;	ram[5123] = 8'h00;
	ram[5124] = 8'h00;	ram[5125] = 8'h00;	ram[5126] = 8'h00;	ram[5127] = 8'h00;
	ram[5128] = 8'h00;	ram[5129] = 8'h00;	ram[5130] = 8'h00;	ram[5131] = 8'h00;
	ram[5132] = 8'h00;	ram[5133] = 8'h00;	ram[5134] = 8'h00;	ram[5135] = 8'h00;
	ram[5136] = 8'h00;	ram[5137] = 8'h00;	ram[5138] = 8'h00;	ram[5139] = 8'h00;
	ram[5140] = 8'h00;	ram[5141] = 8'h00;	ram[5142] = 8'h00;	ram[5143] = 8'h00;
	ram[5144] = 8'h00;	ram[5145] = 8'h00;	ram[5146] = 8'h00;	ram[5147] = 8'h00;
	ram[5148] = 8'h00;	ram[5149] = 8'h00;	ram[5150] = 8'h00;	ram[5151] = 8'h00;
	ram[5152] = 8'h00;	ram[5153] = 8'h00;	ram[5154] = 8'h00;	ram[5155] = 8'h00;
	ram[5156] = 8'h00;	ram[5157] = 8'h00;	ram[5158] = 8'h00;	ram[5159] = 8'h00;
	ram[5160] = 8'h00;	ram[5161] = 8'h00;	ram[5162] = 8'h00;	ram[5163] = 8'h00;
	ram[5164] = 8'h00;	ram[5165] = 8'h00;	ram[5166] = 8'h00;	ram[5167] = 8'h00;
	ram[5168] = 8'h00;	ram[5169] = 8'h00;	ram[5170] = 8'h00;	ram[5171] = 8'h00;
	ram[5172] = 8'h00;	ram[5173] = 8'h00;	ram[5174] = 8'h00;	ram[5175] = 8'h00;
	ram[5176] = 8'h00;	ram[5177] = 8'h00;	ram[5178] = 8'h00;	ram[5179] = 8'h00;
	ram[5180] = 8'h00;	ram[5181] = 8'h00;	ram[5182] = 8'h00;	ram[5183] = 8'h00;
	ram[5184] = 8'h00;	ram[5185] = 8'h00;	ram[5186] = 8'h00;	ram[5187] = 8'h00;
	ram[5188] = 8'h00;	ram[5189] = 8'h00;	ram[5190] = 8'h00;	ram[5191] = 8'h00;
	ram[5192] = 8'h00;	ram[5193] = 8'h00;	ram[5194] = 8'h00;	ram[5195] = 8'h00;
	ram[5196] = 8'h00;	ram[5197] = 8'h00;	ram[5198] = 8'h00;	ram[5199] = 8'h00;
	ram[5200] = 8'h00;	ram[5201] = 8'h00;	ram[5202] = 8'h00;	ram[5203] = 8'h00;
	ram[5204] = 8'h00;	ram[5205] = 8'h00;	ram[5206] = 8'h00;	ram[5207] = 8'h00;
	ram[5208] = 8'h00;	ram[5209] = 8'h00;	ram[5210] = 8'h00;	ram[5211] = 8'h00;
	ram[5212] = 8'h00;	ram[5213] = 8'h00;	ram[5214] = 8'h00;	ram[5215] = 8'h00;
	ram[5216] = 8'h00;	ram[5217] = 8'h00;	ram[5218] = 8'h00;	ram[5219] = 8'h00;
	ram[5220] = 8'h00;	ram[5221] = 8'h00;	ram[5222] = 8'h00;	ram[5223] = 8'h00;
	ram[5224] = 8'h00;	ram[5225] = 8'h00;	ram[5226] = 8'h00;	ram[5227] = 8'h00;
	ram[5228] = 8'h00;	ram[5229] = 8'h00;	ram[5230] = 8'h00;	ram[5231] = 8'h00;
	ram[5232] = 8'h00;	ram[5233] = 8'h00;	ram[5234] = 8'h00;	ram[5235] = 8'h00;
	ram[5236] = 8'h00;	ram[5237] = 8'h00;	ram[5238] = 8'h00;	ram[5239] = 8'h00;
	ram[5240] = 8'h00;	ram[5241] = 8'h00;	ram[5242] = 8'h00;	ram[5243] = 8'h00;
	ram[5244] = 8'h00;	ram[5245] = 8'h00;	ram[5246] = 8'h00;	ram[5247] = 8'h00;
	ram[5248] = 8'h00;	ram[5249] = 8'h00;	ram[5250] = 8'h00;	ram[5251] = 8'h00;
	ram[5252] = 8'h00;	ram[5253] = 8'h00;	ram[5254] = 8'h00;	ram[5255] = 8'h00;
	ram[5256] = 8'h00;	ram[5257] = 8'h00;	ram[5258] = 8'h00;	ram[5259] = 8'h00;
	ram[5260] = 8'h00;	ram[5261] = 8'h00;	ram[5262] = 8'h00;	ram[5263] = 8'h00;
	ram[5264] = 8'h00;	ram[5265] = 8'h00;	ram[5266] = 8'h00;	ram[5267] = 8'h00;
	ram[5268] = 8'h00;	ram[5269] = 8'h00;	ram[5270] = 8'h00;	ram[5271] = 8'h00;
	ram[5272] = 8'h00;	ram[5273] = 8'h00;	ram[5274] = 8'h00;	ram[5275] = 8'h00;
	ram[5276] = 8'h00;	ram[5277] = 8'h00;	ram[5278] = 8'h00;	ram[5279] = 8'h00;
	ram[5280] = 8'h00;	ram[5281] = 8'h00;	ram[5282] = 8'h00;	ram[5283] = 8'h00;
	ram[5284] = 8'h00;	ram[5285] = 8'h00;	ram[5286] = 8'h00;	ram[5287] = 8'h00;
	ram[5288] = 8'h00;	ram[5289] = 8'h00;	ram[5290] = 8'h00;	ram[5291] = 8'h00;
	ram[5292] = 8'h00;	ram[5293] = 8'h00;	ram[5294] = 8'h00;	ram[5295] = 8'h00;
	ram[5296] = 8'h00;	ram[5297] = 8'h00;	ram[5298] = 8'h00;	ram[5299] = 8'h00;
	ram[5300] = 8'h00;	ram[5301] = 8'h00;	ram[5302] = 8'h00;	ram[5303] = 8'h00;
	ram[5304] = 8'h00;	ram[5305] = 8'h00;	ram[5306] = 8'h00;	ram[5307] = 8'h00;
	ram[5308] = 8'h00;	ram[5309] = 8'h00;	ram[5310] = 8'h00;	ram[5311] = 8'h00;
	ram[5312] = 8'h00;	ram[5313] = 8'h00;	ram[5314] = 8'h00;	ram[5315] = 8'h00;
	ram[5316] = 8'h00;	ram[5317] = 8'h00;	ram[5318] = 8'h00;	ram[5319] = 8'h00;
	ram[5320] = 8'h00;	ram[5321] = 8'h00;	ram[5322] = 8'h00;	ram[5323] = 8'h00;
	ram[5324] = 8'h00;	ram[5325] = 8'h00;	ram[5326] = 8'h00;	ram[5327] = 8'h00;
	ram[5328] = 8'h00;	ram[5329] = 8'h00;	ram[5330] = 8'h00;	ram[5331] = 8'h00;
	ram[5332] = 8'h00;	ram[5333] = 8'h00;	ram[5334] = 8'h00;	ram[5335] = 8'h00;
	ram[5336] = 8'h00;	ram[5337] = 8'h00;	ram[5338] = 8'h00;	ram[5339] = 8'h00;
	ram[5340] = 8'h00;	ram[5341] = 8'h00;	ram[5342] = 8'h00;	ram[5343] = 8'h00;
	ram[5344] = 8'h00;	ram[5345] = 8'h00;	ram[5346] = 8'h00;	ram[5347] = 8'h00;
	ram[5348] = 8'h00;	ram[5349] = 8'h00;	ram[5350] = 8'h00;	ram[5351] = 8'h00;
	ram[5352] = 8'h00;	ram[5353] = 8'h00;	ram[5354] = 8'h00;	ram[5355] = 8'h00;
	ram[5356] = 8'h00;	ram[5357] = 8'h00;	ram[5358] = 8'h00;	ram[5359] = 8'h00;
	ram[5360] = 8'h00;	ram[5361] = 8'h00;	ram[5362] = 8'h00;	ram[5363] = 8'h00;
	ram[5364] = 8'h00;	ram[5365] = 8'h00;	ram[5366] = 8'h00;	ram[5367] = 8'h00;
	ram[5368] = 8'h00;	ram[5369] = 8'h00;	ram[5370] = 8'h00;	ram[5371] = 8'h00;
	ram[5372] = 8'h00;	ram[5373] = 8'h00;	ram[5374] = 8'h00;	ram[5375] = 8'h00;
	ram[5376] = 8'h00;	ram[5377] = 8'h00;	ram[5378] = 8'h00;	ram[5379] = 8'h00;
	ram[5380] = 8'h00;	ram[5381] = 8'h00;	ram[5382] = 8'h00;	ram[5383] = 8'h00;
	ram[5384] = 8'h00;	ram[5385] = 8'h00;	ram[5386] = 8'h00;	ram[5387] = 8'h00;
	ram[5388] = 8'h00;	ram[5389] = 8'h00;	ram[5390] = 8'h00;	ram[5391] = 8'h00;
	ram[5392] = 8'h00;	ram[5393] = 8'h00;	ram[5394] = 8'h00;	ram[5395] = 8'h00;
	ram[5396] = 8'h00;	ram[5397] = 8'h00;	ram[5398] = 8'h00;	ram[5399] = 8'h00;
	ram[5400] = 8'h00;	ram[5401] = 8'h00;	ram[5402] = 8'h00;	ram[5403] = 8'h00;
	ram[5404] = 8'h00;	ram[5405] = 8'h00;	ram[5406] = 8'h00;	ram[5407] = 8'h00;
	ram[5408] = 8'h00;	ram[5409] = 8'h00;	ram[5410] = 8'h00;	ram[5411] = 8'h00;
	ram[5412] = 8'h00;	ram[5413] = 8'h00;	ram[5414] = 8'h00;	ram[5415] = 8'h00;
	ram[5416] = 8'h00;	ram[5417] = 8'h00;	ram[5418] = 8'h00;	ram[5419] = 8'h00;
	ram[5420] = 8'h00;	ram[5421] = 8'h00;	ram[5422] = 8'h00;	ram[5423] = 8'h00;
	ram[5424] = 8'h00;	ram[5425] = 8'h00;	ram[5426] = 8'h00;	ram[5427] = 8'h00;
	ram[5428] = 8'h00;	ram[5429] = 8'h00;	ram[5430] = 8'h00;	ram[5431] = 8'h00;
	ram[5432] = 8'h00;	ram[5433] = 8'h00;	ram[5434] = 8'h00;	ram[5435] = 8'h00;
	ram[5436] = 8'h00;	ram[5437] = 8'h00;	ram[5438] = 8'h00;	ram[5439] = 8'h00;
	ram[5440] = 8'h00;	ram[5441] = 8'h00;	ram[5442] = 8'h00;	ram[5443] = 8'h00;
	ram[5444] = 8'h00;	ram[5445] = 8'h00;	ram[5446] = 8'h00;	ram[5447] = 8'h00;
	ram[5448] = 8'h00;	ram[5449] = 8'h00;	ram[5450] = 8'h00;	ram[5451] = 8'h00;
	ram[5452] = 8'h00;	ram[5453] = 8'h00;	ram[5454] = 8'h00;	ram[5455] = 8'h00;
	ram[5456] = 8'h00;	ram[5457] = 8'h00;	ram[5458] = 8'h00;	ram[5459] = 8'h00;
	ram[5460] = 8'h00;	ram[5461] = 8'h00;	ram[5462] = 8'h00;	ram[5463] = 8'h00;
	ram[5464] = 8'h00;	ram[5465] = 8'h00;	ram[5466] = 8'h00;	ram[5467] = 8'h00;
	ram[5468] = 8'h00;	ram[5469] = 8'h00;	ram[5470] = 8'h00;	ram[5471] = 8'h00;
	ram[5472] = 8'h00;	ram[5473] = 8'h00;	ram[5474] = 8'h00;	ram[5475] = 8'h00;
	ram[5476] = 8'h00;	ram[5477] = 8'h00;	ram[5478] = 8'h00;	ram[5479] = 8'h00;
	ram[5480] = 8'h00;	ram[5481] = 8'h00;	ram[5482] = 8'h00;	ram[5483] = 8'h00;
	ram[5484] = 8'h00;	ram[5485] = 8'h00;	ram[5486] = 8'h00;	ram[5487] = 8'h00;
	ram[5488] = 8'h00;	ram[5489] = 8'h00;	ram[5490] = 8'h00;	ram[5491] = 8'h00;
	ram[5492] = 8'h00;	ram[5493] = 8'h00;	ram[5494] = 8'h00;	ram[5495] = 8'h00;
	ram[5496] = 8'h00;	ram[5497] = 8'h00;	ram[5498] = 8'h00;	ram[5499] = 8'h00;
	ram[5500] = 8'h00;	ram[5501] = 8'h00;	ram[5502] = 8'h00;	ram[5503] = 8'h00;
	ram[5504] = 8'h00;	ram[5505] = 8'h00;	ram[5506] = 8'h00;	ram[5507] = 8'h00;
	ram[5508] = 8'h00;	ram[5509] = 8'h00;	ram[5510] = 8'h00;	ram[5511] = 8'h00;
	ram[5512] = 8'h00;	ram[5513] = 8'h00;	ram[5514] = 8'h00;	ram[5515] = 8'h00;
	ram[5516] = 8'h00;	ram[5517] = 8'h00;	ram[5518] = 8'h00;	ram[5519] = 8'h00;
	ram[5520] = 8'h00;	ram[5521] = 8'h00;	ram[5522] = 8'h00;	ram[5523] = 8'h00;
	ram[5524] = 8'h00;	ram[5525] = 8'h00;	ram[5526] = 8'h00;	ram[5527] = 8'h00;
	ram[5528] = 8'h00;	ram[5529] = 8'h00;	ram[5530] = 8'h00;	ram[5531] = 8'h00;
	ram[5532] = 8'h00;	ram[5533] = 8'h00;	ram[5534] = 8'h00;	ram[5535] = 8'h00;
	ram[5536] = 8'h00;	ram[5537] = 8'h00;	ram[5538] = 8'h00;	ram[5539] = 8'h00;
	ram[5540] = 8'h00;	ram[5541] = 8'h00;	ram[5542] = 8'h00;	ram[5543] = 8'h00;
	ram[5544] = 8'h00;	ram[5545] = 8'h00;	ram[5546] = 8'h00;	ram[5547] = 8'h00;
	ram[5548] = 8'h00;	ram[5549] = 8'h00;	ram[5550] = 8'h00;	ram[5551] = 8'h00;
	ram[5552] = 8'h00;	ram[5553] = 8'h00;	ram[5554] = 8'h00;	ram[5555] = 8'h00;
	ram[5556] = 8'h00;	ram[5557] = 8'h00;	ram[5558] = 8'h00;	ram[5559] = 8'h00;
	ram[5560] = 8'h00;	ram[5561] = 8'h00;	ram[5562] = 8'h00;	ram[5563] = 8'h00;
	ram[5564] = 8'h00;	ram[5565] = 8'h00;	ram[5566] = 8'h00;	ram[5567] = 8'h00;
	ram[5568] = 8'h00;	ram[5569] = 8'h00;	ram[5570] = 8'h00;	ram[5571] = 8'h00;
	ram[5572] = 8'h00;	ram[5573] = 8'h00;	ram[5574] = 8'h00;	ram[5575] = 8'h00;
	ram[5576] = 8'h00;	ram[5577] = 8'h00;	ram[5578] = 8'h00;	ram[5579] = 8'h00;
	ram[5580] = 8'h00;	ram[5581] = 8'h00;	ram[5582] = 8'h00;	ram[5583] = 8'h00;
	ram[5584] = 8'h00;	ram[5585] = 8'h00;	ram[5586] = 8'h00;	ram[5587] = 8'h00;
	ram[5588] = 8'h00;	ram[5589] = 8'h00;	ram[5590] = 8'h00;	ram[5591] = 8'h00;
	ram[5592] = 8'h00;	ram[5593] = 8'h00;	ram[5594] = 8'h00;	ram[5595] = 8'h00;
	ram[5596] = 8'h00;	ram[5597] = 8'h00;	ram[5598] = 8'h00;	ram[5599] = 8'h00;
	ram[5600] = 8'h00;	ram[5601] = 8'h00;	ram[5602] = 8'h00;	ram[5603] = 8'h00;
	ram[5604] = 8'h00;	ram[5605] = 8'h00;	ram[5606] = 8'h00;	ram[5607] = 8'h00;
	ram[5608] = 8'h00;	ram[5609] = 8'h00;	ram[5610] = 8'h00;	ram[5611] = 8'h00;
	ram[5612] = 8'h00;	ram[5613] = 8'h00;	ram[5614] = 8'h00;	ram[5615] = 8'h00;
	ram[5616] = 8'h00;	ram[5617] = 8'h00;	ram[5618] = 8'h00;	ram[5619] = 8'h00;
	ram[5620] = 8'h00;	ram[5621] = 8'h00;	ram[5622] = 8'h00;	ram[5623] = 8'h00;
	ram[5624] = 8'h00;	ram[5625] = 8'h00;	ram[5626] = 8'h00;	ram[5627] = 8'h00;
	ram[5628] = 8'h00;	ram[5629] = 8'h00;	ram[5630] = 8'h00;	ram[5631] = 8'h00;
	ram[5632] = 8'h00;	ram[5633] = 8'h00;	ram[5634] = 8'h00;	ram[5635] = 8'h00;
	ram[5636] = 8'h00;	ram[5637] = 8'h00;	ram[5638] = 8'h00;	ram[5639] = 8'h00;
	ram[5640] = 8'h00;	ram[5641] = 8'h00;	ram[5642] = 8'h00;	ram[5643] = 8'h00;
	ram[5644] = 8'h00;	ram[5645] = 8'h00;	ram[5646] = 8'h00;	ram[5647] = 8'h00;
	ram[5648] = 8'h00;	ram[5649] = 8'h00;	ram[5650] = 8'h00;	ram[5651] = 8'h00;
	ram[5652] = 8'h00;	ram[5653] = 8'h00;	ram[5654] = 8'h00;	ram[5655] = 8'h00;
	ram[5656] = 8'h00;	ram[5657] = 8'h00;	ram[5658] = 8'h00;	ram[5659] = 8'h00;
	ram[5660] = 8'h00;	ram[5661] = 8'h00;	ram[5662] = 8'h00;	ram[5663] = 8'h00;
	ram[5664] = 8'h00;	ram[5665] = 8'h00;	ram[5666] = 8'h00;	ram[5667] = 8'h00;
	ram[5668] = 8'h00;	ram[5669] = 8'h00;	ram[5670] = 8'h00;	ram[5671] = 8'h00;
	ram[5672] = 8'h00;	ram[5673] = 8'h00;	ram[5674] = 8'h00;	ram[5675] = 8'h00;
	ram[5676] = 8'h00;	ram[5677] = 8'h00;	ram[5678] = 8'h00;	ram[5679] = 8'h00;
	ram[5680] = 8'h00;	ram[5681] = 8'h00;	ram[5682] = 8'h00;	ram[5683] = 8'h00;
	ram[5684] = 8'h00;	ram[5685] = 8'h00;	ram[5686] = 8'h00;	ram[5687] = 8'h00;
	ram[5688] = 8'h00;	ram[5689] = 8'h00;	ram[5690] = 8'h00;	ram[5691] = 8'h00;
	ram[5692] = 8'h00;	ram[5693] = 8'h00;	ram[5694] = 8'h00;	ram[5695] = 8'h00;
	ram[5696] = 8'h00;	ram[5697] = 8'h00;	ram[5698] = 8'h00;	ram[5699] = 8'h00;
	ram[5700] = 8'h00;	ram[5701] = 8'h00;	ram[5702] = 8'h00;	ram[5703] = 8'h00;
	ram[5704] = 8'h00;	ram[5705] = 8'h00;	ram[5706] = 8'h00;	ram[5707] = 8'h00;
	ram[5708] = 8'h00;	ram[5709] = 8'h00;	ram[5710] = 8'h00;	ram[5711] = 8'h00;
	ram[5712] = 8'h00;	ram[5713] = 8'h00;	ram[5714] = 8'h00;	ram[5715] = 8'h00;
	ram[5716] = 8'h00;	ram[5717] = 8'h00;	ram[5718] = 8'h00;	ram[5719] = 8'h00;
	ram[5720] = 8'h00;	ram[5721] = 8'h00;	ram[5722] = 8'h00;	ram[5723] = 8'h00;
	ram[5724] = 8'h00;	ram[5725] = 8'h00;	ram[5726] = 8'h00;	ram[5727] = 8'h00;
	ram[5728] = 8'h00;	ram[5729] = 8'h00;	ram[5730] = 8'h00;	ram[5731] = 8'h00;
	ram[5732] = 8'h00;	ram[5733] = 8'h00;	ram[5734] = 8'h00;	ram[5735] = 8'h00;
	ram[5736] = 8'h00;	ram[5737] = 8'h00;	ram[5738] = 8'h00;	ram[5739] = 8'h00;
	ram[5740] = 8'h00;	ram[5741] = 8'h00;	ram[5742] = 8'h00;	ram[5743] = 8'h00;
	ram[5744] = 8'h00;	ram[5745] = 8'h00;	ram[5746] = 8'h00;	ram[5747] = 8'h00;
	ram[5748] = 8'h00;	ram[5749] = 8'h00;	ram[5750] = 8'h00;	ram[5751] = 8'h00;
	ram[5752] = 8'h00;	ram[5753] = 8'h00;	ram[5754] = 8'h00;	ram[5755] = 8'h00;
	ram[5756] = 8'h00;	ram[5757] = 8'h00;	ram[5758] = 8'h00;	ram[5759] = 8'h00;
	ram[5760] = 8'h00;	ram[5761] = 8'h00;	ram[5762] = 8'h00;	ram[5763] = 8'h00;
	ram[5764] = 8'h00;	ram[5765] = 8'h00;	ram[5766] = 8'h00;	ram[5767] = 8'h00;
	ram[5768] = 8'h00;	ram[5769] = 8'h00;	ram[5770] = 8'h00;	ram[5771] = 8'h00;
	ram[5772] = 8'h00;	ram[5773] = 8'h00;	ram[5774] = 8'h00;	ram[5775] = 8'h00;
	ram[5776] = 8'h00;	ram[5777] = 8'h00;	ram[5778] = 8'h00;	ram[5779] = 8'h00;
	ram[5780] = 8'h00;	ram[5781] = 8'h00;	ram[5782] = 8'h00;	ram[5783] = 8'h00;
	ram[5784] = 8'h00;	ram[5785] = 8'h00;	ram[5786] = 8'h00;	ram[5787] = 8'h00;
	ram[5788] = 8'h00;	ram[5789] = 8'h00;	ram[5790] = 8'h00;	ram[5791] = 8'h00;
	ram[5792] = 8'h00;	ram[5793] = 8'h00;	ram[5794] = 8'h00;	ram[5795] = 8'h00;
	ram[5796] = 8'h00;	ram[5797] = 8'h00;	ram[5798] = 8'h00;	ram[5799] = 8'h00;
	ram[5800] = 8'h00;	ram[5801] = 8'h00;	ram[5802] = 8'h00;	ram[5803] = 8'h00;
	ram[5804] = 8'h00;	ram[5805] = 8'h00;	ram[5806] = 8'h00;	ram[5807] = 8'h00;
	ram[5808] = 8'h00;	ram[5809] = 8'h00;	ram[5810] = 8'h00;	ram[5811] = 8'h00;
	ram[5812] = 8'h00;	ram[5813] = 8'h00;	ram[5814] = 8'h00;	ram[5815] = 8'h00;
	ram[5816] = 8'h00;	ram[5817] = 8'h00;	ram[5818] = 8'h00;	ram[5819] = 8'h00;
	ram[5820] = 8'h00;	ram[5821] = 8'h00;	ram[5822] = 8'h00;	ram[5823] = 8'h00;
	ram[5824] = 8'h00;	ram[5825] = 8'h00;	ram[5826] = 8'h00;	ram[5827] = 8'h00;
	ram[5828] = 8'h00;	ram[5829] = 8'h00;	ram[5830] = 8'h00;	ram[5831] = 8'h00;
	ram[5832] = 8'h00;	ram[5833] = 8'h00;	ram[5834] = 8'h00;	ram[5835] = 8'h00;
	ram[5836] = 8'h00;	ram[5837] = 8'h00;	ram[5838] = 8'h00;	ram[5839] = 8'h00;
	ram[5840] = 8'h00;	ram[5841] = 8'h00;	ram[5842] = 8'h00;	ram[5843] = 8'h00;
	ram[5844] = 8'h00;	ram[5845] = 8'h00;	ram[5846] = 8'h00;	ram[5847] = 8'h00;
	ram[5848] = 8'h00;	ram[5849] = 8'h00;	ram[5850] = 8'h00;	ram[5851] = 8'h00;
	ram[5852] = 8'h00;	ram[5853] = 8'h00;	ram[5854] = 8'h00;	ram[5855] = 8'h00;
	ram[5856] = 8'h00;	ram[5857] = 8'h00;	ram[5858] = 8'h00;	ram[5859] = 8'h00;
	ram[5860] = 8'h00;	ram[5861] = 8'h00;	ram[5862] = 8'h00;	ram[5863] = 8'h00;
	ram[5864] = 8'h00;	ram[5865] = 8'h00;	ram[5866] = 8'h00;	ram[5867] = 8'h00;
	ram[5868] = 8'h00;	ram[5869] = 8'h00;	ram[5870] = 8'h00;	ram[5871] = 8'h00;
	ram[5872] = 8'h00;	ram[5873] = 8'h00;	ram[5874] = 8'h00;	ram[5875] = 8'h00;
	ram[5876] = 8'h00;	ram[5877] = 8'h00;	ram[5878] = 8'h00;	ram[5879] = 8'h00;
	ram[5880] = 8'h00;	ram[5881] = 8'h00;	ram[5882] = 8'h00;	ram[5883] = 8'h00;
	ram[5884] = 8'h00;	ram[5885] = 8'h00;	ram[5886] = 8'h00;	ram[5887] = 8'h00;
	ram[5888] = 8'h00;	ram[5889] = 8'h00;	ram[5890] = 8'h00;	ram[5891] = 8'h00;
	ram[5892] = 8'h00;	ram[5893] = 8'h00;	ram[5894] = 8'h00;	ram[5895] = 8'h00;
	ram[5896] = 8'h00;	ram[5897] = 8'h00;	ram[5898] = 8'h00;	ram[5899] = 8'h00;
	ram[5900] = 8'h00;	ram[5901] = 8'h00;	ram[5902] = 8'h00;	ram[5903] = 8'h00;
	ram[5904] = 8'h00;	ram[5905] = 8'h00;	ram[5906] = 8'h00;	ram[5907] = 8'h00;
	ram[5908] = 8'h00;	ram[5909] = 8'h00;	ram[5910] = 8'h00;	ram[5911] = 8'h00;
	ram[5912] = 8'h00;	ram[5913] = 8'h00;	ram[5914] = 8'h00;	ram[5915] = 8'h00;
	ram[5916] = 8'h00;	ram[5917] = 8'h00;	ram[5918] = 8'h00;	ram[5919] = 8'h00;
	ram[5920] = 8'h00;	ram[5921] = 8'h00;	ram[5922] = 8'h00;	ram[5923] = 8'h00;
	ram[5924] = 8'h00;	ram[5925] = 8'h00;	ram[5926] = 8'h00;	ram[5927] = 8'h00;
	ram[5928] = 8'h00;	ram[5929] = 8'h00;	ram[5930] = 8'h00;	ram[5931] = 8'h00;
	ram[5932] = 8'h00;	ram[5933] = 8'h00;	ram[5934] = 8'h00;	ram[5935] = 8'h00;
	ram[5936] = 8'h00;	ram[5937] = 8'h00;	ram[5938] = 8'h00;	ram[5939] = 8'h00;
	ram[5940] = 8'h00;	ram[5941] = 8'h00;	ram[5942] = 8'h00;	ram[5943] = 8'h00;
	ram[5944] = 8'h00;	ram[5945] = 8'h00;	ram[5946] = 8'h00;	ram[5947] = 8'h00;
	ram[5948] = 8'h00;	ram[5949] = 8'h00;	ram[5950] = 8'h00;	ram[5951] = 8'h00;
	ram[5952] = 8'h00;	ram[5953] = 8'h00;	ram[5954] = 8'h00;	ram[5955] = 8'h00;
	ram[5956] = 8'h00;	ram[5957] = 8'h00;	ram[5958] = 8'h00;	ram[5959] = 8'h00;
	ram[5960] = 8'h00;	ram[5961] = 8'h00;	ram[5962] = 8'h00;	ram[5963] = 8'h00;
	ram[5964] = 8'h00;	ram[5965] = 8'h00;	ram[5966] = 8'h00;	ram[5967] = 8'h00;
	ram[5968] = 8'h00;	ram[5969] = 8'h00;	ram[5970] = 8'h00;	ram[5971] = 8'h00;
	ram[5972] = 8'h00;	ram[5973] = 8'h00;	ram[5974] = 8'h00;	ram[5975] = 8'h00;
	ram[5976] = 8'h00;	ram[5977] = 8'h00;	ram[5978] = 8'h00;	ram[5979] = 8'h00;
	ram[5980] = 8'h00;	ram[5981] = 8'h00;	ram[5982] = 8'h00;	ram[5983] = 8'h00;
	ram[5984] = 8'h00;	ram[5985] = 8'h00;	ram[5986] = 8'h00;	ram[5987] = 8'h00;
	ram[5988] = 8'h00;	ram[5989] = 8'h00;	ram[5990] = 8'h00;	ram[5991] = 8'h00;
	ram[5992] = 8'h00;	ram[5993] = 8'h00;	ram[5994] = 8'h00;	ram[5995] = 8'h00;
	ram[5996] = 8'h00;	ram[5997] = 8'h00;	ram[5998] = 8'h00;	ram[5999] = 8'h00;
	ram[6000] = 8'h00;	ram[6001] = 8'h00;	ram[6002] = 8'h00;	ram[6003] = 8'h00;
	ram[6004] = 8'h00;	ram[6005] = 8'h00;	ram[6006] = 8'h00;	ram[6007] = 8'h00;
	ram[6008] = 8'h00;	ram[6009] = 8'h00;	ram[6010] = 8'h00;	ram[6011] = 8'h00;
	ram[6012] = 8'h00;	ram[6013] = 8'h00;	ram[6014] = 8'h00;	ram[6015] = 8'h00;
	ram[6016] = 8'h00;	ram[6017] = 8'h00;	ram[6018] = 8'h00;	ram[6019] = 8'h00;
	ram[6020] = 8'h00;	ram[6021] = 8'h00;	ram[6022] = 8'h00;	ram[6023] = 8'h00;
	ram[6024] = 8'h00;	ram[6025] = 8'h00;	ram[6026] = 8'h00;	ram[6027] = 8'h00;
	ram[6028] = 8'h00;	ram[6029] = 8'h00;	ram[6030] = 8'h00;	ram[6031] = 8'h00;
	ram[6032] = 8'h00;	ram[6033] = 8'h00;	ram[6034] = 8'h00;	ram[6035] = 8'h00;
	ram[6036] = 8'h00;	ram[6037] = 8'h00;	ram[6038] = 8'h00;	ram[6039] = 8'h00;
	ram[6040] = 8'h00;	ram[6041] = 8'h00;	ram[6042] = 8'h00;	ram[6043] = 8'h00;
	ram[6044] = 8'h00;	ram[6045] = 8'h00;	ram[6046] = 8'h00;	ram[6047] = 8'h00;
	ram[6048] = 8'h00;	ram[6049] = 8'h00;	ram[6050] = 8'h00;	ram[6051] = 8'h00;
	ram[6052] = 8'h00;	ram[6053] = 8'h00;	ram[6054] = 8'h00;	ram[6055] = 8'h00;
	ram[6056] = 8'h00;	ram[6057] = 8'h00;	ram[6058] = 8'h00;	ram[6059] = 8'h00;
	ram[6060] = 8'h00;	ram[6061] = 8'h00;	ram[6062] = 8'h00;	ram[6063] = 8'h00;
	ram[6064] = 8'h00;	ram[6065] = 8'h00;	ram[6066] = 8'h00;	ram[6067] = 8'h00;
	ram[6068] = 8'h00;	ram[6069] = 8'h00;	ram[6070] = 8'h00;	ram[6071] = 8'h00;
	ram[6072] = 8'h00;	ram[6073] = 8'h00;	ram[6074] = 8'h00;	ram[6075] = 8'h00;
	ram[6076] = 8'h00;	ram[6077] = 8'h00;	ram[6078] = 8'h00;	ram[6079] = 8'h00;
	ram[6080] = 8'h00;	ram[6081] = 8'h00;	ram[6082] = 8'h00;	ram[6083] = 8'h00;
	ram[6084] = 8'h00;	ram[6085] = 8'h00;	ram[6086] = 8'h00;	ram[6087] = 8'h00;
	ram[6088] = 8'h00;	ram[6089] = 8'h00;	ram[6090] = 8'h00;	ram[6091] = 8'h00;
	ram[6092] = 8'h00;	ram[6093] = 8'h00;	ram[6094] = 8'h00;	ram[6095] = 8'h00;
	ram[6096] = 8'h00;	ram[6097] = 8'h00;	ram[6098] = 8'h00;	ram[6099] = 8'h00;
	ram[6100] = 8'h00;	ram[6101] = 8'h00;	ram[6102] = 8'h00;	ram[6103] = 8'h00;
	ram[6104] = 8'h00;	ram[6105] = 8'h00;	ram[6106] = 8'h00;	ram[6107] = 8'h00;
	ram[6108] = 8'h00;	ram[6109] = 8'h00;	ram[6110] = 8'h00;	ram[6111] = 8'h00;
	ram[6112] = 8'h00;	ram[6113] = 8'h00;	ram[6114] = 8'h00;	ram[6115] = 8'h00;
	ram[6116] = 8'h00;	ram[6117] = 8'h00;	ram[6118] = 8'h00;	ram[6119] = 8'h00;
	ram[6120] = 8'h00;	ram[6121] = 8'h00;	ram[6122] = 8'h00;	ram[6123] = 8'h00;
	ram[6124] = 8'h00;	ram[6125] = 8'h00;	ram[6126] = 8'h00;	ram[6127] = 8'h00;
	ram[6128] = 8'h00;	ram[6129] = 8'h00;	ram[6130] = 8'h00;	ram[6131] = 8'h00;
	ram[6132] = 8'h00;	ram[6133] = 8'h00;	ram[6134] = 8'h00;	ram[6135] = 8'h00;
	ram[6136] = 8'h00;	ram[6137] = 8'h00;	ram[6138] = 8'h00;	ram[6139] = 8'h00;
	ram[6140] = 8'h00;	ram[6141] = 8'h00;	ram[6142] = 8'h00;	ram[6143] = 8'h00;
	ram[6144] = 8'h00;	ram[6145] = 8'h00;	ram[6146] = 8'h00;	ram[6147] = 8'h00;
	ram[6148] = 8'h00;	ram[6149] = 8'h00;	ram[6150] = 8'h00;	ram[6151] = 8'h00;
	ram[6152] = 8'h00;	ram[6153] = 8'h00;	ram[6154] = 8'h00;	ram[6155] = 8'h00;
	ram[6156] = 8'h00;	ram[6157] = 8'h00;	ram[6158] = 8'h00;	ram[6159] = 8'h00;
	ram[6160] = 8'h00;	ram[6161] = 8'h00;	ram[6162] = 8'h00;	ram[6163] = 8'h00;
	ram[6164] = 8'h00;	ram[6165] = 8'h00;	ram[6166] = 8'h00;	ram[6167] = 8'h00;
	ram[6168] = 8'h00;	ram[6169] = 8'h00;	ram[6170] = 8'h00;	ram[6171] = 8'h00;
	ram[6172] = 8'h00;	ram[6173] = 8'h00;	ram[6174] = 8'h00;	ram[6175] = 8'h00;
	ram[6176] = 8'h00;	ram[6177] = 8'h00;	ram[6178] = 8'h00;	ram[6179] = 8'h00;
	ram[6180] = 8'h00;	ram[6181] = 8'h00;	ram[6182] = 8'h00;	ram[6183] = 8'h00;
	ram[6184] = 8'h00;	ram[6185] = 8'h00;	ram[6186] = 8'h00;	ram[6187] = 8'h00;
	ram[6188] = 8'h00;	ram[6189] = 8'h00;	ram[6190] = 8'h00;	ram[6191] = 8'h00;
	ram[6192] = 8'h00;	ram[6193] = 8'h00;	ram[6194] = 8'h00;	ram[6195] = 8'h00;
	ram[6196] = 8'h00;	ram[6197] = 8'h00;	ram[6198] = 8'h00;	ram[6199] = 8'h00;
	ram[6200] = 8'h00;	ram[6201] = 8'h00;	ram[6202] = 8'h00;	ram[6203] = 8'h00;
	ram[6204] = 8'h00;	ram[6205] = 8'h00;	ram[6206] = 8'h00;	ram[6207] = 8'h00;
	ram[6208] = 8'h00;	ram[6209] = 8'h00;	ram[6210] = 8'h00;	ram[6211] = 8'h00;
	ram[6212] = 8'h00;	ram[6213] = 8'h00;	ram[6214] = 8'h00;	ram[6215] = 8'h00;
	ram[6216] = 8'h00;	ram[6217] = 8'h00;	ram[6218] = 8'h00;	ram[6219] = 8'h00;
	ram[6220] = 8'h00;	ram[6221] = 8'h00;	ram[6222] = 8'h00;	ram[6223] = 8'h00;
	ram[6224] = 8'h00;	ram[6225] = 8'h00;	ram[6226] = 8'h00;	ram[6227] = 8'h00;
	ram[6228] = 8'h00;	ram[6229] = 8'h00;	ram[6230] = 8'h00;	ram[6231] = 8'h00;
	ram[6232] = 8'h00;	ram[6233] = 8'h00;	ram[6234] = 8'h00;	ram[6235] = 8'h00;
	ram[6236] = 8'h00;	ram[6237] = 8'h00;	ram[6238] = 8'h00;	ram[6239] = 8'h00;
	ram[6240] = 8'h00;	ram[6241] = 8'h00;	ram[6242] = 8'h00;	ram[6243] = 8'h00;
	ram[6244] = 8'h00;	ram[6245] = 8'h00;	ram[6246] = 8'h00;	ram[6247] = 8'h00;
	ram[6248] = 8'h00;	ram[6249] = 8'h00;	ram[6250] = 8'h00;	ram[6251] = 8'h00;
	ram[6252] = 8'h00;	ram[6253] = 8'h00;	ram[6254] = 8'h00;	ram[6255] = 8'h00;
	ram[6256] = 8'h00;	ram[6257] = 8'h00;	ram[6258] = 8'h00;	ram[6259] = 8'h00;
	ram[6260] = 8'h00;	ram[6261] = 8'h00;	ram[6262] = 8'h00;	ram[6263] = 8'h00;
	ram[6264] = 8'h00;	ram[6265] = 8'h00;	ram[6266] = 8'h00;	ram[6267] = 8'h00;
	ram[6268] = 8'h00;	ram[6269] = 8'h00;	ram[6270] = 8'h00;	ram[6271] = 8'h00;
	ram[6272] = 8'h00;	ram[6273] = 8'h00;	ram[6274] = 8'h00;	ram[6275] = 8'h00;
	ram[6276] = 8'h00;	ram[6277] = 8'h00;	ram[6278] = 8'h00;	ram[6279] = 8'h00;
	ram[6280] = 8'h00;	ram[6281] = 8'h00;	ram[6282] = 8'h00;	ram[6283] = 8'h00;
	ram[6284] = 8'h00;	ram[6285] = 8'h00;	ram[6286] = 8'h00;	ram[6287] = 8'h00;
	ram[6288] = 8'h00;	ram[6289] = 8'h00;	ram[6290] = 8'h00;	ram[6291] = 8'h00;
	ram[6292] = 8'h00;	ram[6293] = 8'h00;	ram[6294] = 8'h00;	ram[6295] = 8'h00;
	ram[6296] = 8'h00;	ram[6297] = 8'h00;	ram[6298] = 8'h00;	ram[6299] = 8'h00;
	ram[6300] = 8'h00;	ram[6301] = 8'h00;	ram[6302] = 8'h00;	ram[6303] = 8'h00;
	ram[6304] = 8'h00;	ram[6305] = 8'h00;	ram[6306] = 8'h00;	ram[6307] = 8'h00;
	ram[6308] = 8'h00;	ram[6309] = 8'h00;	ram[6310] = 8'h00;	ram[6311] = 8'h00;
	ram[6312] = 8'h00;	ram[6313] = 8'h00;	ram[6314] = 8'h00;	ram[6315] = 8'h00;
	ram[6316] = 8'h00;	ram[6317] = 8'h00;	ram[6318] = 8'h00;	ram[6319] = 8'h00;
	ram[6320] = 8'h00;	ram[6321] = 8'h00;	ram[6322] = 8'h00;	ram[6323] = 8'h00;
	ram[6324] = 8'h00;	ram[6325] = 8'h00;	ram[6326] = 8'h00;	ram[6327] = 8'h00;
	ram[6328] = 8'h00;	ram[6329] = 8'h00;	ram[6330] = 8'h00;	ram[6331] = 8'h00;
	ram[6332] = 8'h00;	ram[6333] = 8'h00;	ram[6334] = 8'h00;	ram[6335] = 8'h00;
	ram[6336] = 8'h00;	ram[6337] = 8'h00;	ram[6338] = 8'h00;	ram[6339] = 8'h00;
	ram[6340] = 8'h00;	ram[6341] = 8'h00;	ram[6342] = 8'h00;	ram[6343] = 8'h00;
	ram[6344] = 8'h00;	ram[6345] = 8'h00;	ram[6346] = 8'h00;	ram[6347] = 8'h00;
	ram[6348] = 8'h00;	ram[6349] = 8'h00;	ram[6350] = 8'h00;	ram[6351] = 8'h00;
	ram[6352] = 8'h00;	ram[6353] = 8'h00;	ram[6354] = 8'h00;	ram[6355] = 8'h00;
	ram[6356] = 8'h00;	ram[6357] = 8'h00;	ram[6358] = 8'h00;	ram[6359] = 8'h00;
	ram[6360] = 8'h00;	ram[6361] = 8'h00;	ram[6362] = 8'h00;	ram[6363] = 8'h00;
	ram[6364] = 8'h00;	ram[6365] = 8'h00;	ram[6366] = 8'h00;	ram[6367] = 8'h00;
	ram[6368] = 8'h00;	ram[6369] = 8'h00;	ram[6370] = 8'h00;	ram[6371] = 8'h00;
	ram[6372] = 8'h00;	ram[6373] = 8'h00;	ram[6374] = 8'h00;	ram[6375] = 8'h00;
	ram[6376] = 8'h00;	ram[6377] = 8'h00;	ram[6378] = 8'h00;	ram[6379] = 8'h00;
	ram[6380] = 8'h00;	ram[6381] = 8'h00;	ram[6382] = 8'h00;	ram[6383] = 8'h00;
	ram[6384] = 8'h00;	ram[6385] = 8'h00;	ram[6386] = 8'h00;	ram[6387] = 8'h00;
	ram[6388] = 8'h00;	ram[6389] = 8'h00;	ram[6390] = 8'h00;	ram[6391] = 8'h00;
	ram[6392] = 8'h00;	ram[6393] = 8'h00;	ram[6394] = 8'h00;	ram[6395] = 8'h00;
	ram[6396] = 8'h00;	ram[6397] = 8'h00;	ram[6398] = 8'h00;	ram[6399] = 8'h00;
	ram[6400] = 8'h00;	ram[6401] = 8'h00;	ram[6402] = 8'h00;	ram[6403] = 8'h00;
	ram[6404] = 8'h00;	ram[6405] = 8'h00;	ram[6406] = 8'h00;	ram[6407] = 8'h00;
	ram[6408] = 8'h00;	ram[6409] = 8'h00;	ram[6410] = 8'h00;	ram[6411] = 8'h00;
	ram[6412] = 8'h00;	ram[6413] = 8'h00;	ram[6414] = 8'h00;	ram[6415] = 8'h00;
	ram[6416] = 8'h00;	ram[6417] = 8'h00;	ram[6418] = 8'h00;	ram[6419] = 8'h00;
	ram[6420] = 8'h00;	ram[6421] = 8'h00;	ram[6422] = 8'h00;	ram[6423] = 8'h00;
	ram[6424] = 8'h00;	ram[6425] = 8'h00;	ram[6426] = 8'h00;	ram[6427] = 8'h00;
	ram[6428] = 8'h00;	ram[6429] = 8'h00;	ram[6430] = 8'h00;	ram[6431] = 8'h00;
	ram[6432] = 8'h00;	ram[6433] = 8'h00;	ram[6434] = 8'h00;	ram[6435] = 8'h00;
	ram[6436] = 8'h00;	ram[6437] = 8'h00;	ram[6438] = 8'h00;	ram[6439] = 8'h00;
	ram[6440] = 8'h00;	ram[6441] = 8'h00;	ram[6442] = 8'h00;	ram[6443] = 8'h00;
	ram[6444] = 8'h00;	ram[6445] = 8'h00;	ram[6446] = 8'h00;	ram[6447] = 8'h00;
	ram[6448] = 8'h00;	ram[6449] = 8'h00;	ram[6450] = 8'h00;	ram[6451] = 8'h00;
	ram[6452] = 8'h00;	ram[6453] = 8'h00;	ram[6454] = 8'h00;	ram[6455] = 8'h00;
	ram[6456] = 8'h00;	ram[6457] = 8'h00;	ram[6458] = 8'h00;	ram[6459] = 8'h00;
	ram[6460] = 8'h00;	ram[6461] = 8'h00;	ram[6462] = 8'h00;	ram[6463] = 8'h00;
	ram[6464] = 8'h00;	ram[6465] = 8'h00;	ram[6466] = 8'h00;	ram[6467] = 8'h00;
	ram[6468] = 8'h00;	ram[6469] = 8'h00;	ram[6470] = 8'h00;	ram[6471] = 8'h00;
	ram[6472] = 8'h00;	ram[6473] = 8'h00;	ram[6474] = 8'h00;	ram[6475] = 8'h00;
	ram[6476] = 8'h00;	ram[6477] = 8'h00;	ram[6478] = 8'h00;	ram[6479] = 8'h00;
	ram[6480] = 8'h00;	ram[6481] = 8'h00;	ram[6482] = 8'h00;	ram[6483] = 8'h00;
	ram[6484] = 8'h00;	ram[6485] = 8'h00;	ram[6486] = 8'h00;	ram[6487] = 8'h00;
	ram[6488] = 8'h00;	ram[6489] = 8'h00;	ram[6490] = 8'h00;	ram[6491] = 8'h00;
	ram[6492] = 8'h00;	ram[6493] = 8'h00;	ram[6494] = 8'h00;	ram[6495] = 8'h00;
	ram[6496] = 8'h00;	ram[6497] = 8'h00;	ram[6498] = 8'h00;	ram[6499] = 8'h00;
	ram[6500] = 8'h00;	ram[6501] = 8'h00;	ram[6502] = 8'h00;	ram[6503] = 8'h00;
	ram[6504] = 8'h00;	ram[6505] = 8'h00;	ram[6506] = 8'h00;	ram[6507] = 8'h00;
	ram[6508] = 8'h00;	ram[6509] = 8'h00;	ram[6510] = 8'h00;	ram[6511] = 8'h00;
	ram[6512] = 8'h00;	ram[6513] = 8'h00;	ram[6514] = 8'h00;	ram[6515] = 8'h00;
	ram[6516] = 8'h00;	ram[6517] = 8'h00;	ram[6518] = 8'h00;	ram[6519] = 8'h00;
	ram[6520] = 8'h00;	ram[6521] = 8'h00;	ram[6522] = 8'h00;	ram[6523] = 8'h00;
	ram[6524] = 8'h00;	ram[6525] = 8'h00;	ram[6526] = 8'h00;	ram[6527] = 8'h00;
	ram[6528] = 8'h00;	ram[6529] = 8'h00;	ram[6530] = 8'h00;	ram[6531] = 8'h00;
	ram[6532] = 8'h00;	ram[6533] = 8'h00;	ram[6534] = 8'h00;	ram[6535] = 8'h00;
	ram[6536] = 8'h00;	ram[6537] = 8'h00;	ram[6538] = 8'h00;	ram[6539] = 8'h00;
	ram[6540] = 8'h00;	ram[6541] = 8'h00;	ram[6542] = 8'h00;	ram[6543] = 8'h00;
	ram[6544] = 8'h00;	ram[6545] = 8'h00;	ram[6546] = 8'h00;	ram[6547] = 8'h00;
	ram[6548] = 8'h00;	ram[6549] = 8'h00;	ram[6550] = 8'h00;	ram[6551] = 8'h00;
	ram[6552] = 8'h00;	ram[6553] = 8'h00;	ram[6554] = 8'h00;	ram[6555] = 8'h00;
	ram[6556] = 8'h00;	ram[6557] = 8'h00;	ram[6558] = 8'h00;	ram[6559] = 8'h00;
	ram[6560] = 8'h00;	ram[6561] = 8'h00;	ram[6562] = 8'h00;	ram[6563] = 8'h00;
	ram[6564] = 8'h00;	ram[6565] = 8'h00;	ram[6566] = 8'h00;	ram[6567] = 8'h00;
	ram[6568] = 8'h00;	ram[6569] = 8'h00;	ram[6570] = 8'h00;	ram[6571] = 8'h00;
	ram[6572] = 8'h00;	ram[6573] = 8'h00;	ram[6574] = 8'h00;	ram[6575] = 8'h00;
	ram[6576] = 8'h00;	ram[6577] = 8'h00;	ram[6578] = 8'h00;	ram[6579] = 8'h00;
	ram[6580] = 8'h00;	ram[6581] = 8'h00;	ram[6582] = 8'h00;	ram[6583] = 8'h00;
	ram[6584] = 8'h00;	ram[6585] = 8'h00;	ram[6586] = 8'h00;	ram[6587] = 8'h00;
	ram[6588] = 8'h00;	ram[6589] = 8'h00;	ram[6590] = 8'h00;	ram[6591] = 8'h00;
	ram[6592] = 8'h00;	ram[6593] = 8'h00;	ram[6594] = 8'h00;	ram[6595] = 8'h00;
	ram[6596] = 8'h00;	ram[6597] = 8'h00;	ram[6598] = 8'h00;	ram[6599] = 8'h00;
	ram[6600] = 8'h00;	ram[6601] = 8'h00;	ram[6602] = 8'h00;	ram[6603] = 8'h00;
	ram[6604] = 8'h00;	ram[6605] = 8'h00;	ram[6606] = 8'h00;	ram[6607] = 8'h00;
	ram[6608] = 8'h00;	ram[6609] = 8'h00;	ram[6610] = 8'h00;	ram[6611] = 8'h00;
	ram[6612] = 8'h00;	ram[6613] = 8'h00;	ram[6614] = 8'h00;	ram[6615] = 8'h00;
	ram[6616] = 8'h00;	ram[6617] = 8'h00;	ram[6618] = 8'h00;	ram[6619] = 8'h00;
	ram[6620] = 8'h00;	ram[6621] = 8'h00;	ram[6622] = 8'h00;	ram[6623] = 8'h00;
	ram[6624] = 8'h00;	ram[6625] = 8'h00;	ram[6626] = 8'h00;	ram[6627] = 8'h00;
	ram[6628] = 8'h00;	ram[6629] = 8'h00;	ram[6630] = 8'h00;	ram[6631] = 8'h00;
	ram[6632] = 8'h00;	ram[6633] = 8'h00;	ram[6634] = 8'h00;	ram[6635] = 8'h00;
	ram[6636] = 8'h00;	ram[6637] = 8'h00;	ram[6638] = 8'h00;	ram[6639] = 8'h00;
	ram[6640] = 8'h00;	ram[6641] = 8'h00;	ram[6642] = 8'h00;	ram[6643] = 8'h00;
	ram[6644] = 8'h00;	ram[6645] = 8'h00;	ram[6646] = 8'h00;	ram[6647] = 8'h00;
	ram[6648] = 8'h00;	ram[6649] = 8'h00;	ram[6650] = 8'h00;	ram[6651] = 8'h00;
	ram[6652] = 8'h00;	ram[6653] = 8'h00;	ram[6654] = 8'h00;	ram[6655] = 8'h00;
	ram[6656] = 8'h00;	ram[6657] = 8'h00;	ram[6658] = 8'h00;	ram[6659] = 8'h00;
	ram[6660] = 8'h00;	ram[6661] = 8'h00;	ram[6662] = 8'h00;	ram[6663] = 8'h00;
	ram[6664] = 8'h00;	ram[6665] = 8'h00;	ram[6666] = 8'h00;	ram[6667] = 8'h00;
	ram[6668] = 8'h00;	ram[6669] = 8'h00;	ram[6670] = 8'h00;	ram[6671] = 8'h00;
	ram[6672] = 8'h00;	ram[6673] = 8'h00;	ram[6674] = 8'h00;	ram[6675] = 8'h00;
	ram[6676] = 8'h00;	ram[6677] = 8'h00;	ram[6678] = 8'h00;	ram[6679] = 8'h00;
	ram[6680] = 8'h00;	ram[6681] = 8'h00;	ram[6682] = 8'h00;	ram[6683] = 8'h00;
	ram[6684] = 8'h00;	ram[6685] = 8'h00;	ram[6686] = 8'h00;	ram[6687] = 8'h00;
	ram[6688] = 8'h00;	ram[6689] = 8'h00;	ram[6690] = 8'h00;	ram[6691] = 8'h00;
	ram[6692] = 8'h00;	ram[6693] = 8'h00;	ram[6694] = 8'h00;	ram[6695] = 8'h00;
	ram[6696] = 8'h00;	ram[6697] = 8'h00;	ram[6698] = 8'h00;	ram[6699] = 8'h00;
	ram[6700] = 8'h00;	ram[6701] = 8'h00;	ram[6702] = 8'h00;	ram[6703] = 8'h00;
	ram[6704] = 8'h00;	ram[6705] = 8'h00;	ram[6706] = 8'h00;	ram[6707] = 8'h00;
	ram[6708] = 8'h00;	ram[6709] = 8'h00;	ram[6710] = 8'h00;	ram[6711] = 8'h00;
	ram[6712] = 8'h00;	ram[6713] = 8'h00;	ram[6714] = 8'h00;	ram[6715] = 8'h00;
	ram[6716] = 8'h00;	ram[6717] = 8'h00;	ram[6718] = 8'h00;	ram[6719] = 8'h00;
	ram[6720] = 8'h00;	ram[6721] = 8'h00;	ram[6722] = 8'h00;	ram[6723] = 8'h00;
	ram[6724] = 8'h00;	ram[6725] = 8'h00;	ram[6726] = 8'h00;	ram[6727] = 8'h00;
	ram[6728] = 8'h00;	ram[6729] = 8'h00;	ram[6730] = 8'h00;	ram[6731] = 8'h00;
	ram[6732] = 8'h00;	ram[6733] = 8'h00;	ram[6734] = 8'h00;	ram[6735] = 8'h00;
	ram[6736] = 8'h00;	ram[6737] = 8'h00;	ram[6738] = 8'h00;	ram[6739] = 8'h00;
	ram[6740] = 8'h00;	ram[6741] = 8'h00;	ram[6742] = 8'h00;	ram[6743] = 8'h00;
	ram[6744] = 8'h00;	ram[6745] = 8'h00;	ram[6746] = 8'h00;	ram[6747] = 8'h00;
	ram[6748] = 8'h00;	ram[6749] = 8'h00;	ram[6750] = 8'h00;	ram[6751] = 8'h00;
	ram[6752] = 8'h00;	ram[6753] = 8'h00;	ram[6754] = 8'h00;	ram[6755] = 8'h00;
	ram[6756] = 8'h00;	ram[6757] = 8'h00;	ram[6758] = 8'h00;	ram[6759] = 8'h00;
	ram[6760] = 8'h00;	ram[6761] = 8'h00;	ram[6762] = 8'h00;	ram[6763] = 8'h00;
	ram[6764] = 8'h00;	ram[6765] = 8'h00;	ram[6766] = 8'h00;	ram[6767] = 8'h00;
	ram[6768] = 8'h00;	ram[6769] = 8'h00;	ram[6770] = 8'h00;	ram[6771] = 8'h00;
	ram[6772] = 8'h00;	ram[6773] = 8'h00;	ram[6774] = 8'h00;	ram[6775] = 8'h00;
	ram[6776] = 8'h00;	ram[6777] = 8'h00;	ram[6778] = 8'h00;	ram[6779] = 8'h00;
	ram[6780] = 8'h00;	ram[6781] = 8'h00;	ram[6782] = 8'h00;	ram[6783] = 8'h00;
	ram[6784] = 8'h00;	ram[6785] = 8'h00;	ram[6786] = 8'h00;	ram[6787] = 8'h00;
	ram[6788] = 8'h00;	ram[6789] = 8'h00;	ram[6790] = 8'h00;	ram[6791] = 8'h00;
	ram[6792] = 8'h00;	ram[6793] = 8'h00;	ram[6794] = 8'h00;	ram[6795] = 8'h00;
	ram[6796] = 8'h00;	ram[6797] = 8'h00;	ram[6798] = 8'h00;	ram[6799] = 8'h00;
	ram[6800] = 8'h00;	ram[6801] = 8'h00;	ram[6802] = 8'h00;	ram[6803] = 8'h00;
	ram[6804] = 8'h00;	ram[6805] = 8'h00;	ram[6806] = 8'h00;	ram[6807] = 8'h00;
	ram[6808] = 8'h00;	ram[6809] = 8'h00;	ram[6810] = 8'h00;	ram[6811] = 8'h00;
	ram[6812] = 8'h00;	ram[6813] = 8'h00;	ram[6814] = 8'h00;	ram[6815] = 8'h00;
	ram[6816] = 8'h00;	ram[6817] = 8'h00;	ram[6818] = 8'h00;	ram[6819] = 8'h00;
	ram[6820] = 8'h00;	ram[6821] = 8'h00;	ram[6822] = 8'h00;	ram[6823] = 8'h00;
	ram[6824] = 8'h00;	ram[6825] = 8'h00;	ram[6826] = 8'h00;	ram[6827] = 8'h00;
	ram[6828] = 8'h00;	ram[6829] = 8'h00;	ram[6830] = 8'h00;	ram[6831] = 8'h00;
	ram[6832] = 8'h00;	ram[6833] = 8'h00;	ram[6834] = 8'h00;	ram[6835] = 8'h00;
	ram[6836] = 8'h00;	ram[6837] = 8'h00;	ram[6838] = 8'h00;	ram[6839] = 8'h00;
	ram[6840] = 8'h00;	ram[6841] = 8'h00;	ram[6842] = 8'h00;	ram[6843] = 8'h00;
	ram[6844] = 8'h00;	ram[6845] = 8'h00;	ram[6846] = 8'h00;	ram[6847] = 8'h00;
	ram[6848] = 8'h00;	ram[6849] = 8'h00;	ram[6850] = 8'h00;	ram[6851] = 8'h00;
	ram[6852] = 8'h00;	ram[6853] = 8'h00;	ram[6854] = 8'h00;	ram[6855] = 8'h00;
	ram[6856] = 8'h00;	ram[6857] = 8'h00;	ram[6858] = 8'h00;	ram[6859] = 8'h00;
	ram[6860] = 8'h00;	ram[6861] = 8'h00;	ram[6862] = 8'h00;	ram[6863] = 8'h00;
	ram[6864] = 8'h00;	ram[6865] = 8'h00;	ram[6866] = 8'h00;	ram[6867] = 8'h00;
	ram[6868] = 8'h00;	ram[6869] = 8'h00;	ram[6870] = 8'h00;	ram[6871] = 8'h00;
	ram[6872] = 8'h00;	ram[6873] = 8'h00;	ram[6874] = 8'h00;	ram[6875] = 8'h00;
	ram[6876] = 8'h00;	ram[6877] = 8'h00;	ram[6878] = 8'h00;	ram[6879] = 8'h00;
	ram[6880] = 8'h00;	ram[6881] = 8'h00;	ram[6882] = 8'h00;	ram[6883] = 8'h00;
	ram[6884] = 8'h00;	ram[6885] = 8'h00;	ram[6886] = 8'h00;	ram[6887] = 8'h00;
	ram[6888] = 8'h00;	ram[6889] = 8'h00;	ram[6890] = 8'h00;	ram[6891] = 8'h00;
	ram[6892] = 8'h00;	ram[6893] = 8'h00;	ram[6894] = 8'h00;	ram[6895] = 8'h00;
	ram[6896] = 8'h00;	ram[6897] = 8'h00;	ram[6898] = 8'h00;	ram[6899] = 8'h00;
	ram[6900] = 8'h00;	ram[6901] = 8'h00;	ram[6902] = 8'h00;	ram[6903] = 8'h00;
	ram[6904] = 8'h00;	ram[6905] = 8'h00;	ram[6906] = 8'h00;	ram[6907] = 8'h00;
	ram[6908] = 8'h00;	ram[6909] = 8'h00;	ram[6910] = 8'h00;	ram[6911] = 8'h00;
	ram[6912] = 8'h00;	ram[6913] = 8'h00;	ram[6914] = 8'h00;	ram[6915] = 8'h00;
	ram[6916] = 8'h00;	ram[6917] = 8'h00;	ram[6918] = 8'h00;	ram[6919] = 8'h00;
	ram[6920] = 8'h00;	ram[6921] = 8'h00;	ram[6922] = 8'h00;	ram[6923] = 8'h00;
	ram[6924] = 8'h00;	ram[6925] = 8'h00;	ram[6926] = 8'h00;	ram[6927] = 8'h00;
	ram[6928] = 8'h00;	ram[6929] = 8'h00;	ram[6930] = 8'h00;	ram[6931] = 8'h00;
	ram[6932] = 8'h00;	ram[6933] = 8'h00;	ram[6934] = 8'h00;	ram[6935] = 8'h00;
	ram[6936] = 8'h00;	ram[6937] = 8'h00;	ram[6938] = 8'h00;	ram[6939] = 8'h00;
	ram[6940] = 8'h00;	ram[6941] = 8'h00;	ram[6942] = 8'h00;	ram[6943] = 8'h00;
	ram[6944] = 8'h00;	ram[6945] = 8'h00;	ram[6946] = 8'h00;	ram[6947] = 8'h00;
	ram[6948] = 8'h00;	ram[6949] = 8'h00;	ram[6950] = 8'h00;	ram[6951] = 8'h00;
	ram[6952] = 8'h00;	ram[6953] = 8'h00;	ram[6954] = 8'h00;	ram[6955] = 8'h00;
	ram[6956] = 8'h00;	ram[6957] = 8'h00;	ram[6958] = 8'h00;	ram[6959] = 8'h00;
	ram[6960] = 8'h00;	ram[6961] = 8'h00;	ram[6962] = 8'h00;	ram[6963] = 8'h00;
	ram[6964] = 8'h00;	ram[6965] = 8'h00;	ram[6966] = 8'h00;	ram[6967] = 8'h00;
	ram[6968] = 8'h00;	ram[6969] = 8'h00;	ram[6970] = 8'h00;	ram[6971] = 8'h00;
	ram[6972] = 8'h00;	ram[6973] = 8'h00;	ram[6974] = 8'h00;	ram[6975] = 8'h00;
	ram[6976] = 8'h00;	ram[6977] = 8'h00;	ram[6978] = 8'h00;	ram[6979] = 8'h00;
	ram[6980] = 8'h00;	ram[6981] = 8'h00;	ram[6982] = 8'h00;	ram[6983] = 8'h00;
	ram[6984] = 8'h00;	ram[6985] = 8'h00;	ram[6986] = 8'h00;	ram[6987] = 8'h00;
	ram[6988] = 8'h00;	ram[6989] = 8'h00;	ram[6990] = 8'h00;	ram[6991] = 8'h00;
	ram[6992] = 8'h00;	ram[6993] = 8'h00;	ram[6994] = 8'h00;	ram[6995] = 8'h00;
	ram[6996] = 8'h00;	ram[6997] = 8'h00;	ram[6998] = 8'h00;	ram[6999] = 8'h00;
	ram[7000] = 8'h00;	ram[7001] = 8'h00;	ram[7002] = 8'h00;	ram[7003] = 8'h00;
	ram[7004] = 8'h00;	ram[7005] = 8'h00;	ram[7006] = 8'h00;	ram[7007] = 8'h00;
	ram[7008] = 8'h00;	ram[7009] = 8'h00;	ram[7010] = 8'h00;	ram[7011] = 8'h00;
	ram[7012] = 8'h00;	ram[7013] = 8'h00;	ram[7014] = 8'h00;	ram[7015] = 8'h00;
	ram[7016] = 8'h00;	ram[7017] = 8'h00;	ram[7018] = 8'h00;	ram[7019] = 8'h00;
	ram[7020] = 8'h00;	ram[7021] = 8'h00;	ram[7022] = 8'h00;	ram[7023] = 8'h00;
	ram[7024] = 8'h00;	ram[7025] = 8'h00;	ram[7026] = 8'h00;	ram[7027] = 8'h00;
	ram[7028] = 8'h00;	ram[7029] = 8'h00;	ram[7030] = 8'h00;	ram[7031] = 8'h00;
	ram[7032] = 8'h00;	ram[7033] = 8'h00;	ram[7034] = 8'h00;	ram[7035] = 8'h00;
	ram[7036] = 8'h00;	ram[7037] = 8'h00;	ram[7038] = 8'h00;	ram[7039] = 8'h00;
	ram[7040] = 8'h00;	ram[7041] = 8'h00;	ram[7042] = 8'h00;	ram[7043] = 8'h00;
	ram[7044] = 8'h00;	ram[7045] = 8'h00;	ram[7046] = 8'h00;	ram[7047] = 8'h00;
	ram[7048] = 8'h00;	ram[7049] = 8'h00;	ram[7050] = 8'h00;	ram[7051] = 8'h00;
	ram[7052] = 8'h00;	ram[7053] = 8'h00;	ram[7054] = 8'h00;	ram[7055] = 8'h00;
	ram[7056] = 8'h00;	ram[7057] = 8'h00;	ram[7058] = 8'h00;	ram[7059] = 8'h00;
	ram[7060] = 8'h00;	ram[7061] = 8'h00;	ram[7062] = 8'h00;	ram[7063] = 8'h00;
	ram[7064] = 8'h00;	ram[7065] = 8'h00;	ram[7066] = 8'h00;	ram[7067] = 8'h00;
	ram[7068] = 8'h00;	ram[7069] = 8'h00;	ram[7070] = 8'h00;	ram[7071] = 8'h00;
	ram[7072] = 8'h00;	ram[7073] = 8'h00;	ram[7074] = 8'h00;	ram[7075] = 8'h00;
	ram[7076] = 8'h00;	ram[7077] = 8'h00;	ram[7078] = 8'h00;	ram[7079] = 8'h00;
	ram[7080] = 8'h00;	ram[7081] = 8'h00;	ram[7082] = 8'h00;	ram[7083] = 8'h00;
	ram[7084] = 8'h00;	ram[7085] = 8'h00;	ram[7086] = 8'h00;	ram[7087] = 8'h00;
	ram[7088] = 8'h00;	ram[7089] = 8'h00;	ram[7090] = 8'h00;	ram[7091] = 8'h00;
	ram[7092] = 8'h00;	ram[7093] = 8'h00;	ram[7094] = 8'h00;	ram[7095] = 8'h00;
	ram[7096] = 8'h00;	ram[7097] = 8'h00;	ram[7098] = 8'h00;	ram[7099] = 8'h00;
	ram[7100] = 8'h00;	ram[7101] = 8'h00;	ram[7102] = 8'h00;	ram[7103] = 8'h00;
	ram[7104] = 8'h00;	ram[7105] = 8'h00;	ram[7106] = 8'h00;	ram[7107] = 8'h00;
	ram[7108] = 8'h00;	ram[7109] = 8'h00;	ram[7110] = 8'h00;	ram[7111] = 8'h00;
	ram[7112] = 8'h00;	ram[7113] = 8'h00;	ram[7114] = 8'h00;	ram[7115] = 8'h00;
	ram[7116] = 8'h00;	ram[7117] = 8'h00;	ram[7118] = 8'h00;	ram[7119] = 8'h00;
	ram[7120] = 8'h00;	ram[7121] = 8'h00;	ram[7122] = 8'h00;	ram[7123] = 8'h00;
	ram[7124] = 8'h00;	ram[7125] = 8'h00;	ram[7126] = 8'h00;	ram[7127] = 8'h00;
	ram[7128] = 8'h00;	ram[7129] = 8'h00;	ram[7130] = 8'h00;	ram[7131] = 8'h00;
	ram[7132] = 8'h00;	ram[7133] = 8'h00;	ram[7134] = 8'h00;	ram[7135] = 8'h00;
	ram[7136] = 8'h00;	ram[7137] = 8'h00;	ram[7138] = 8'h00;	ram[7139] = 8'h00;
	ram[7140] = 8'h00;	ram[7141] = 8'h00;	ram[7142] = 8'h00;	ram[7143] = 8'h00;
	ram[7144] = 8'h00;	ram[7145] = 8'h00;	ram[7146] = 8'h00;	ram[7147] = 8'h00;
	ram[7148] = 8'h00;	ram[7149] = 8'h00;	ram[7150] = 8'h00;	ram[7151] = 8'h00;
	ram[7152] = 8'h00;	ram[7153] = 8'h00;	ram[7154] = 8'h00;	ram[7155] = 8'h00;
	ram[7156] = 8'h00;	ram[7157] = 8'h00;	ram[7158] = 8'h00;	ram[7159] = 8'h00;
	ram[7160] = 8'h00;	ram[7161] = 8'h00;	ram[7162] = 8'h00;	ram[7163] = 8'h00;
	ram[7164] = 8'h00;	ram[7165] = 8'h00;	ram[7166] = 8'h00;	ram[7167] = 8'h00;
	ram[7168] = 8'h00;	ram[7169] = 8'h00;	ram[7170] = 8'h00;	ram[7171] = 8'h00;
	ram[7172] = 8'h00;	ram[7173] = 8'h00;	ram[7174] = 8'h00;	ram[7175] = 8'h00;
	ram[7176] = 8'h00;	ram[7177] = 8'h00;	ram[7178] = 8'h00;	ram[7179] = 8'h00;
	ram[7180] = 8'h00;	ram[7181] = 8'h00;	ram[7182] = 8'h00;	ram[7183] = 8'h00;
	ram[7184] = 8'h00;	ram[7185] = 8'h00;	ram[7186] = 8'h00;	ram[7187] = 8'h00;
	ram[7188] = 8'h00;	ram[7189] = 8'h00;	ram[7190] = 8'h00;	ram[7191] = 8'h00;
	ram[7192] = 8'h00;	ram[7193] = 8'h00;	ram[7194] = 8'h00;	ram[7195] = 8'h00;
	ram[7196] = 8'h00;	ram[7197] = 8'h00;	ram[7198] = 8'h00;	ram[7199] = 8'h00;
	ram[7200] = 8'h00;	ram[7201] = 8'h00;	ram[7202] = 8'h00;	ram[7203] = 8'h00;
	ram[7204] = 8'h00;	ram[7205] = 8'h00;	ram[7206] = 8'h00;	ram[7207] = 8'h00;
	ram[7208] = 8'h00;	ram[7209] = 8'h00;	ram[7210] = 8'h00;	ram[7211] = 8'h00;
	ram[7212] = 8'h00;	ram[7213] = 8'h00;	ram[7214] = 8'h00;	ram[7215] = 8'h00;
	ram[7216] = 8'h00;	ram[7217] = 8'h00;	ram[7218] = 8'h00;	ram[7219] = 8'h00;
	ram[7220] = 8'h00;	ram[7221] = 8'h00;	ram[7222] = 8'h00;	ram[7223] = 8'h00;
	ram[7224] = 8'h00;	ram[7225] = 8'h00;	ram[7226] = 8'h00;	ram[7227] = 8'h00;
	ram[7228] = 8'h00;	ram[7229] = 8'h00;	ram[7230] = 8'h00;	ram[7231] = 8'h00;
	ram[7232] = 8'h00;	ram[7233] = 8'h00;	ram[7234] = 8'h00;	ram[7235] = 8'h00;
	ram[7236] = 8'h00;	ram[7237] = 8'h00;	ram[7238] = 8'h00;	ram[7239] = 8'h00;
	ram[7240] = 8'h00;	ram[7241] = 8'h00;	ram[7242] = 8'h00;	ram[7243] = 8'h00;
	ram[7244] = 8'h00;	ram[7245] = 8'h00;	ram[7246] = 8'h00;	ram[7247] = 8'h00;
	ram[7248] = 8'h00;	ram[7249] = 8'h00;	ram[7250] = 8'h00;	ram[7251] = 8'h00;
	ram[7252] = 8'h00;	ram[7253] = 8'h00;	ram[7254] = 8'h00;	ram[7255] = 8'h00;
	ram[7256] = 8'h00;	ram[7257] = 8'h00;	ram[7258] = 8'h00;	ram[7259] = 8'h00;
	ram[7260] = 8'h00;	ram[7261] = 8'h00;	ram[7262] = 8'h00;	ram[7263] = 8'h00;
	ram[7264] = 8'h00;	ram[7265] = 8'h00;	ram[7266] = 8'h00;	ram[7267] = 8'h00;
	ram[7268] = 8'h00;	ram[7269] = 8'h00;	ram[7270] = 8'h00;	ram[7271] = 8'h00;
	ram[7272] = 8'h00;	ram[7273] = 8'h00;	ram[7274] = 8'h00;	ram[7275] = 8'h00;
	ram[7276] = 8'h00;	ram[7277] = 8'h00;	ram[7278] = 8'h00;	ram[7279] = 8'h00;
	ram[7280] = 8'h00;	ram[7281] = 8'h00;	ram[7282] = 8'h00;	ram[7283] = 8'h00;
	ram[7284] = 8'h00;	ram[7285] = 8'h00;	ram[7286] = 8'h00;	ram[7287] = 8'h00;
	ram[7288] = 8'h00;	ram[7289] = 8'h00;	ram[7290] = 8'h00;	ram[7291] = 8'h00;
	ram[7292] = 8'h00;	ram[7293] = 8'h00;	ram[7294] = 8'h00;	ram[7295] = 8'h00;
	ram[7296] = 8'h00;	ram[7297] = 8'h00;	ram[7298] = 8'h00;	ram[7299] = 8'h00;
	ram[7300] = 8'h00;	ram[7301] = 8'h00;	ram[7302] = 8'h00;	ram[7303] = 8'h00;
	ram[7304] = 8'h00;	ram[7305] = 8'h00;	ram[7306] = 8'h00;	ram[7307] = 8'h00;
	ram[7308] = 8'h00;	ram[7309] = 8'h00;	ram[7310] = 8'h00;	ram[7311] = 8'h00;
	ram[7312] = 8'h00;	ram[7313] = 8'h00;	ram[7314] = 8'h00;	ram[7315] = 8'h00;
	ram[7316] = 8'h00;	ram[7317] = 8'h00;	ram[7318] = 8'h00;	ram[7319] = 8'h00;
	ram[7320] = 8'h00;	ram[7321] = 8'h00;	ram[7322] = 8'h00;	ram[7323] = 8'h00;
	ram[7324] = 8'h00;	ram[7325] = 8'h00;	ram[7326] = 8'h00;	ram[7327] = 8'h00;
	ram[7328] = 8'h00;	ram[7329] = 8'h00;	ram[7330] = 8'h00;	ram[7331] = 8'h00;
	ram[7332] = 8'h00;	ram[7333] = 8'h00;	ram[7334] = 8'h00;	ram[7335] = 8'h00;
	ram[7336] = 8'h00;	ram[7337] = 8'h00;	ram[7338] = 8'h00;	ram[7339] = 8'h00;
	ram[7340] = 8'h00;	ram[7341] = 8'h00;	ram[7342] = 8'h00;	ram[7343] = 8'h00;
	ram[7344] = 8'h00;	ram[7345] = 8'h00;	ram[7346] = 8'h00;	ram[7347] = 8'h00;
	ram[7348] = 8'h00;	ram[7349] = 8'h00;	ram[7350] = 8'h00;	ram[7351] = 8'h00;
	ram[7352] = 8'h00;	ram[7353] = 8'h00;	ram[7354] = 8'h00;	ram[7355] = 8'h00;
	ram[7356] = 8'h00;	ram[7357] = 8'h00;	ram[7358] = 8'h00;	ram[7359] = 8'h00;
	ram[7360] = 8'h00;	ram[7361] = 8'h00;	ram[7362] = 8'h00;	ram[7363] = 8'h00;
	ram[7364] = 8'h00;	ram[7365] = 8'h00;	ram[7366] = 8'h00;	ram[7367] = 8'h00;
	ram[7368] = 8'h00;	ram[7369] = 8'h00;	ram[7370] = 8'h00;	ram[7371] = 8'h00;
	ram[7372] = 8'h00;	ram[7373] = 8'h00;	ram[7374] = 8'h00;	ram[7375] = 8'h00;
	ram[7376] = 8'h00;	ram[7377] = 8'h00;	ram[7378] = 8'h00;	ram[7379] = 8'h00;
	ram[7380] = 8'h00;	ram[7381] = 8'h00;	ram[7382] = 8'h00;	ram[7383] = 8'h00;
	ram[7384] = 8'h00;	ram[7385] = 8'h00;	ram[7386] = 8'h00;	ram[7387] = 8'h00;
	ram[7388] = 8'h00;	ram[7389] = 8'h00;	ram[7390] = 8'h00;	ram[7391] = 8'h00;
	ram[7392] = 8'h00;	ram[7393] = 8'h00;	ram[7394] = 8'h00;	ram[7395] = 8'h00;
	ram[7396] = 8'h00;	ram[7397] = 8'h00;	ram[7398] = 8'h00;	ram[7399] = 8'h00;
	ram[7400] = 8'h00;	ram[7401] = 8'h00;	ram[7402] = 8'h00;	ram[7403] = 8'h00;
	ram[7404] = 8'h00;	ram[7405] = 8'h00;	ram[7406] = 8'h00;	ram[7407] = 8'h00;
	ram[7408] = 8'h00;	ram[7409] = 8'h00;	ram[7410] = 8'h00;	ram[7411] = 8'h00;
	ram[7412] = 8'h00;	ram[7413] = 8'h00;	ram[7414] = 8'h00;	ram[7415] = 8'h00;
	ram[7416] = 8'h00;	ram[7417] = 8'h00;	ram[7418] = 8'h00;	ram[7419] = 8'h00;
	ram[7420] = 8'h00;	ram[7421] = 8'h00;	ram[7422] = 8'h00;	ram[7423] = 8'h00;
	ram[7424] = 8'h00;	ram[7425] = 8'h00;	ram[7426] = 8'h00;	ram[7427] = 8'h00;
	ram[7428] = 8'h00;	ram[7429] = 8'h00;	ram[7430] = 8'h00;	ram[7431] = 8'h00;
	ram[7432] = 8'h00;	ram[7433] = 8'h00;	ram[7434] = 8'h00;	ram[7435] = 8'h00;
	ram[7436] = 8'h00;	ram[7437] = 8'h00;	ram[7438] = 8'h00;	ram[7439] = 8'h00;
	ram[7440] = 8'h00;	ram[7441] = 8'h00;	ram[7442] = 8'h00;	ram[7443] = 8'h00;
	ram[7444] = 8'h00;	ram[7445] = 8'h00;	ram[7446] = 8'h00;	ram[7447] = 8'h00;
	ram[7448] = 8'h00;	ram[7449] = 8'h00;	ram[7450] = 8'h00;	ram[7451] = 8'h00;
	ram[7452] = 8'h00;	ram[7453] = 8'h00;	ram[7454] = 8'h00;	ram[7455] = 8'h00;
	ram[7456] = 8'h00;	ram[7457] = 8'h00;	ram[7458] = 8'h00;	ram[7459] = 8'h00;
	ram[7460] = 8'h00;	ram[7461] = 8'h00;	ram[7462] = 8'h00;	ram[7463] = 8'h00;
	ram[7464] = 8'h00;	ram[7465] = 8'h00;	ram[7466] = 8'h00;	ram[7467] = 8'h00;
	ram[7468] = 8'h00;	ram[7469] = 8'h00;	ram[7470] = 8'h00;	ram[7471] = 8'h00;
	ram[7472] = 8'h00;	ram[7473] = 8'h00;	ram[7474] = 8'h00;	ram[7475] = 8'h00;
	ram[7476] = 8'h00;	ram[7477] = 8'h00;	ram[7478] = 8'h00;	ram[7479] = 8'h00;
	ram[7480] = 8'h00;	ram[7481] = 8'h00;	ram[7482] = 8'h00;	ram[7483] = 8'h00;
	ram[7484] = 8'h00;	ram[7485] = 8'h00;	ram[7486] = 8'h00;	ram[7487] = 8'h00;
	ram[7488] = 8'h00;	ram[7489] = 8'h00;	ram[7490] = 8'h00;	ram[7491] = 8'h00;
	ram[7492] = 8'h00;	ram[7493] = 8'h00;	ram[7494] = 8'h00;	ram[7495] = 8'h00;
	ram[7496] = 8'h00;	ram[7497] = 8'h00;	ram[7498] = 8'h00;	ram[7499] = 8'h00;
	ram[7500] = 8'h00;	ram[7501] = 8'h00;	ram[7502] = 8'h00;	ram[7503] = 8'h00;
	ram[7504] = 8'h00;	ram[7505] = 8'h00;	ram[7506] = 8'h00;	ram[7507] = 8'h00;
	ram[7508] = 8'h00;	ram[7509] = 8'h00;	ram[7510] = 8'h00;	ram[7511] = 8'h00;
	ram[7512] = 8'h00;	ram[7513] = 8'h00;	ram[7514] = 8'h00;	ram[7515] = 8'h00;
	ram[7516] = 8'h00;	ram[7517] = 8'h00;	ram[7518] = 8'h00;	ram[7519] = 8'h00;
	ram[7520] = 8'h00;	ram[7521] = 8'h00;	ram[7522] = 8'h00;	ram[7523] = 8'h00;
	ram[7524] = 8'h00;	ram[7525] = 8'h00;	ram[7526] = 8'h00;	ram[7527] = 8'h00;
	ram[7528] = 8'h00;	ram[7529] = 8'h00;	ram[7530] = 8'h00;	ram[7531] = 8'h00;
	ram[7532] = 8'h00;	ram[7533] = 8'h00;	ram[7534] = 8'h00;	ram[7535] = 8'h00;
	ram[7536] = 8'h00;	ram[7537] = 8'h00;	ram[7538] = 8'h00;	ram[7539] = 8'h00;
	ram[7540] = 8'h00;	ram[7541] = 8'h00;	ram[7542] = 8'h00;	ram[7543] = 8'h00;
	ram[7544] = 8'h00;	ram[7545] = 8'h00;	ram[7546] = 8'h00;	ram[7547] = 8'h00;
	ram[7548] = 8'h00;	ram[7549] = 8'h00;	ram[7550] = 8'h00;	ram[7551] = 8'h00;
	ram[7552] = 8'h00;	ram[7553] = 8'h00;	ram[7554] = 8'h00;	ram[7555] = 8'h00;
	ram[7556] = 8'h00;	ram[7557] = 8'h00;	ram[7558] = 8'h00;	ram[7559] = 8'h00;
	ram[7560] = 8'h00;	ram[7561] = 8'h00;	ram[7562] = 8'h00;	ram[7563] = 8'h00;
	ram[7564] = 8'h00;	ram[7565] = 8'h00;	ram[7566] = 8'h00;	ram[7567] = 8'h00;
	ram[7568] = 8'h00;	ram[7569] = 8'h00;	ram[7570] = 8'h00;	ram[7571] = 8'h00;
	ram[7572] = 8'h00;	ram[7573] = 8'h00;	ram[7574] = 8'h00;	ram[7575] = 8'h00;
	ram[7576] = 8'h00;	ram[7577] = 8'h00;	ram[7578] = 8'h00;	ram[7579] = 8'h00;
	ram[7580] = 8'h00;	ram[7581] = 8'h00;	ram[7582] = 8'h00;	ram[7583] = 8'h00;
	ram[7584] = 8'h00;	ram[7585] = 8'h00;	ram[7586] = 8'h00;	ram[7587] = 8'h00;
	ram[7588] = 8'h00;	ram[7589] = 8'h00;	ram[7590] = 8'h00;	ram[7591] = 8'h00;
	ram[7592] = 8'h00;	ram[7593] = 8'h00;	ram[7594] = 8'h00;	ram[7595] = 8'h00;
	ram[7596] = 8'h00;	ram[7597] = 8'h00;	ram[7598] = 8'h00;	ram[7599] = 8'h00;
	ram[7600] = 8'h00;	ram[7601] = 8'h00;	ram[7602] = 8'h00;	ram[7603] = 8'h00;
	ram[7604] = 8'h00;	ram[7605] = 8'h00;	ram[7606] = 8'h00;	ram[7607] = 8'h00;
	ram[7608] = 8'h00;	ram[7609] = 8'h00;	ram[7610] = 8'h00;	ram[7611] = 8'h00;
	ram[7612] = 8'h00;	ram[7613] = 8'h00;	ram[7614] = 8'h00;	ram[7615] = 8'h00;
	ram[7616] = 8'h00;	ram[7617] = 8'h00;	ram[7618] = 8'h00;	ram[7619] = 8'h00;
	ram[7620] = 8'h00;	ram[7621] = 8'h00;	ram[7622] = 8'h00;	ram[7623] = 8'h00;
	ram[7624] = 8'h00;	ram[7625] = 8'h00;	ram[7626] = 8'h00;	ram[7627] = 8'h00;
	ram[7628] = 8'h00;	ram[7629] = 8'h00;	ram[7630] = 8'h00;	ram[7631] = 8'h00;
	ram[7632] = 8'h00;	ram[7633] = 8'h00;	ram[7634] = 8'h00;	ram[7635] = 8'h00;
	ram[7636] = 8'h00;	ram[7637] = 8'h00;	ram[7638] = 8'h00;	ram[7639] = 8'h00;
	ram[7640] = 8'h00;	ram[7641] = 8'h00;	ram[7642] = 8'h00;	ram[7643] = 8'h00;
	ram[7644] = 8'h00;	ram[7645] = 8'h00;	ram[7646] = 8'h00;	ram[7647] = 8'h00;
	ram[7648] = 8'h00;	ram[7649] = 8'h00;	ram[7650] = 8'h00;	ram[7651] = 8'h00;
	ram[7652] = 8'h00;	ram[7653] = 8'h00;	ram[7654] = 8'h00;	ram[7655] = 8'h00;
	ram[7656] = 8'h00;	ram[7657] = 8'h00;	ram[7658] = 8'h00;	ram[7659] = 8'h00;
	ram[7660] = 8'h00;	ram[7661] = 8'h00;	ram[7662] = 8'h00;	ram[7663] = 8'h00;
	ram[7664] = 8'h00;	ram[7665] = 8'h00;	ram[7666] = 8'h00;	ram[7667] = 8'h00;
	ram[7668] = 8'h00;	ram[7669] = 8'h00;	ram[7670] = 8'h00;	ram[7671] = 8'h00;
	ram[7672] = 8'h00;	ram[7673] = 8'h00;	ram[7674] = 8'h00;	ram[7675] = 8'h00;
	ram[7676] = 8'h00;	ram[7677] = 8'h00;	ram[7678] = 8'h00;	ram[7679] = 8'h00;
	ram[7680] = 8'h00;	ram[7681] = 8'h00;	ram[7682] = 8'h00;	ram[7683] = 8'h00;
	ram[7684] = 8'h00;	ram[7685] = 8'h00;	ram[7686] = 8'h00;	ram[7687] = 8'h00;
	ram[7688] = 8'h00;	ram[7689] = 8'h00;	ram[7690] = 8'h00;	ram[7691] = 8'h00;
	ram[7692] = 8'h00;	ram[7693] = 8'h00;	ram[7694] = 8'h00;	ram[7695] = 8'h00;
	ram[7696] = 8'h00;	ram[7697] = 8'h00;	ram[7698] = 8'h00;	ram[7699] = 8'h00;
	ram[7700] = 8'h00;	ram[7701] = 8'h00;	ram[7702] = 8'h00;	ram[7703] = 8'h00;
	ram[7704] = 8'h00;	ram[7705] = 8'h00;	ram[7706] = 8'h00;	ram[7707] = 8'h00;
	ram[7708] = 8'h00;	ram[7709] = 8'h00;	ram[7710] = 8'h00;	ram[7711] = 8'h00;
	ram[7712] = 8'h00;	ram[7713] = 8'h00;	ram[7714] = 8'h00;	ram[7715] = 8'h00;
	ram[7716] = 8'h00;	ram[7717] = 8'h00;	ram[7718] = 8'h00;	ram[7719] = 8'h00;
	ram[7720] = 8'h00;	ram[7721] = 8'h00;	ram[7722] = 8'h00;	ram[7723] = 8'h00;
	ram[7724] = 8'h00;	ram[7725] = 8'h00;	ram[7726] = 8'h00;	ram[7727] = 8'h00;
	ram[7728] = 8'h00;	ram[7729] = 8'h00;	ram[7730] = 8'h00;	ram[7731] = 8'h00;
	ram[7732] = 8'h00;	ram[7733] = 8'h00;	ram[7734] = 8'h00;	ram[7735] = 8'h00;
	ram[7736] = 8'h00;	ram[7737] = 8'h00;	ram[7738] = 8'h00;	ram[7739] = 8'h00;
	ram[7740] = 8'h00;	ram[7741] = 8'h00;	ram[7742] = 8'h00;	ram[7743] = 8'h00;
	ram[7744] = 8'h00;	ram[7745] = 8'h00;	ram[7746] = 8'h00;	ram[7747] = 8'h00;
	ram[7748] = 8'h00;	ram[7749] = 8'h00;	ram[7750] = 8'h00;	ram[7751] = 8'h00;
	ram[7752] = 8'h00;	ram[7753] = 8'h00;	ram[7754] = 8'h00;	ram[7755] = 8'h00;
	ram[7756] = 8'h00;	ram[7757] = 8'h00;	ram[7758] = 8'h00;	ram[7759] = 8'h00;
	ram[7760] = 8'h00;	ram[7761] = 8'h00;	ram[7762] = 8'h00;	ram[7763] = 8'h00;
	ram[7764] = 8'h00;	ram[7765] = 8'h00;	ram[7766] = 8'h00;	ram[7767] = 8'h00;
	ram[7768] = 8'h00;	ram[7769] = 8'h00;	ram[7770] = 8'h00;	ram[7771] = 8'h00;
	ram[7772] = 8'h00;	ram[7773] = 8'h00;	ram[7774] = 8'h00;	ram[7775] = 8'h00;
	ram[7776] = 8'h00;	ram[7777] = 8'h00;	ram[7778] = 8'h00;	ram[7779] = 8'h00;
	ram[7780] = 8'h00;	ram[7781] = 8'h00;	ram[7782] = 8'h00;	ram[7783] = 8'h00;
	ram[7784] = 8'h00;	ram[7785] = 8'h00;	ram[7786] = 8'h00;	ram[7787] = 8'h00;
	ram[7788] = 8'h00;	ram[7789] = 8'h00;	ram[7790] = 8'h00;	ram[7791] = 8'h00;
	ram[7792] = 8'h00;	ram[7793] = 8'h00;	ram[7794] = 8'h00;	ram[7795] = 8'h00;
	ram[7796] = 8'h00;	ram[7797] = 8'h00;	ram[7798] = 8'h00;	ram[7799] = 8'h00;
	ram[7800] = 8'h00;	ram[7801] = 8'h00;	ram[7802] = 8'h00;	ram[7803] = 8'h00;
	ram[7804] = 8'h00;	ram[7805] = 8'h00;	ram[7806] = 8'h00;	ram[7807] = 8'h00;
	ram[7808] = 8'h00;	ram[7809] = 8'h00;	ram[7810] = 8'h00;	ram[7811] = 8'h00;
	ram[7812] = 8'h00;	ram[7813] = 8'h00;	ram[7814] = 8'h00;	ram[7815] = 8'h00;
	ram[7816] = 8'h00;	ram[7817] = 8'h00;	ram[7818] = 8'h00;	ram[7819] = 8'h00;
	ram[7820] = 8'h00;	ram[7821] = 8'h00;	ram[7822] = 8'h00;	ram[7823] = 8'h00;
	ram[7824] = 8'h00;	ram[7825] = 8'h00;	ram[7826] = 8'h00;	ram[7827] = 8'h00;
	ram[7828] = 8'h00;	ram[7829] = 8'h00;	ram[7830] = 8'h00;	ram[7831] = 8'h00;
	ram[7832] = 8'h00;	ram[7833] = 8'h00;	ram[7834] = 8'h00;	ram[7835] = 8'h00;
	ram[7836] = 8'h00;	ram[7837] = 8'h00;	ram[7838] = 8'h00;	ram[7839] = 8'h00;
	ram[7840] = 8'h00;	ram[7841] = 8'h00;	ram[7842] = 8'h00;	ram[7843] = 8'h00;
	ram[7844] = 8'h00;	ram[7845] = 8'h00;	ram[7846] = 8'h00;	ram[7847] = 8'h00;
	ram[7848] = 8'h00;	ram[7849] = 8'h00;	ram[7850] = 8'h00;	ram[7851] = 8'h00;
	ram[7852] = 8'h00;	ram[7853] = 8'h00;	ram[7854] = 8'h00;	ram[7855] = 8'h00;
	ram[7856] = 8'h00;	ram[7857] = 8'h00;	ram[7858] = 8'h00;	ram[7859] = 8'h00;
	ram[7860] = 8'h00;	ram[7861] = 8'h00;	ram[7862] = 8'h00;	ram[7863] = 8'h00;
	ram[7864] = 8'h00;	ram[7865] = 8'h00;	ram[7866] = 8'h00;	ram[7867] = 8'h00;
	ram[7868] = 8'h00;	ram[7869] = 8'h00;	ram[7870] = 8'h00;	ram[7871] = 8'h00;
	ram[7872] = 8'h00;	ram[7873] = 8'h00;	ram[7874] = 8'h00;	ram[7875] = 8'h00;
	ram[7876] = 8'h00;	ram[7877] = 8'h00;	ram[7878] = 8'h00;	ram[7879] = 8'h00;
	ram[7880] = 8'h00;	ram[7881] = 8'h00;	ram[7882] = 8'h00;	ram[7883] = 8'h00;
	ram[7884] = 8'h00;	ram[7885] = 8'h00;	ram[7886] = 8'h00;	ram[7887] = 8'h00;
	ram[7888] = 8'h00;	ram[7889] = 8'h00;	ram[7890] = 8'h00;	ram[7891] = 8'h00;
	ram[7892] = 8'h00;	ram[7893] = 8'h00;	ram[7894] = 8'h00;	ram[7895] = 8'h00;
	ram[7896] = 8'h00;	ram[7897] = 8'h00;	ram[7898] = 8'h00;	ram[7899] = 8'h00;
	ram[7900] = 8'h00;	ram[7901] = 8'h00;	ram[7902] = 8'h00;	ram[7903] = 8'h00;
	ram[7904] = 8'h00;	ram[7905] = 8'h00;	ram[7906] = 8'h00;	ram[7907] = 8'h00;
	ram[7908] = 8'h00;	ram[7909] = 8'h00;	ram[7910] = 8'h00;	ram[7911] = 8'h00;
	ram[7912] = 8'h00;	ram[7913] = 8'h00;	ram[7914] = 8'h00;	ram[7915] = 8'h00;
	ram[7916] = 8'h00;	ram[7917] = 8'h00;	ram[7918] = 8'h00;	ram[7919] = 8'h00;
	ram[7920] = 8'h00;	ram[7921] = 8'h00;	ram[7922] = 8'h00;	ram[7923] = 8'h00;
	ram[7924] = 8'h00;	ram[7925] = 8'h00;	ram[7926] = 8'h00;	ram[7927] = 8'h00;
	ram[7928] = 8'h00;	ram[7929] = 8'h00;	ram[7930] = 8'h00;	ram[7931] = 8'h00;
	ram[7932] = 8'h00;	ram[7933] = 8'h00;	ram[7934] = 8'h00;	ram[7935] = 8'h00;
	ram[7936] = 8'h00;	ram[7937] = 8'h00;	ram[7938] = 8'h00;	ram[7939] = 8'h00;
	ram[7940] = 8'h00;	ram[7941] = 8'h00;	ram[7942] = 8'h00;	ram[7943] = 8'h00;
	ram[7944] = 8'h00;	ram[7945] = 8'h00;	ram[7946] = 8'h00;	ram[7947] = 8'h00;
	ram[7948] = 8'h00;	ram[7949] = 8'h00;	ram[7950] = 8'h00;	ram[7951] = 8'h00;
	ram[7952] = 8'h00;	ram[7953] = 8'h00;	ram[7954] = 8'h00;	ram[7955] = 8'h00;
	ram[7956] = 8'h00;	ram[7957] = 8'h00;	ram[7958] = 8'h00;	ram[7959] = 8'h00;
	ram[7960] = 8'h00;	ram[7961] = 8'h00;	ram[7962] = 8'h00;	ram[7963] = 8'h00;
	ram[7964] = 8'h00;	ram[7965] = 8'h00;	ram[7966] = 8'h00;	ram[7967] = 8'h00;
	ram[7968] = 8'h00;	ram[7969] = 8'h00;	ram[7970] = 8'h00;	ram[7971] = 8'h00;
	ram[7972] = 8'h00;	ram[7973] = 8'h00;	ram[7974] = 8'h00;	ram[7975] = 8'h00;
	ram[7976] = 8'h00;	ram[7977] = 8'h00;	ram[7978] = 8'h00;	ram[7979] = 8'h00;
	ram[7980] = 8'h00;	ram[7981] = 8'h00;	ram[7982] = 8'h00;	ram[7983] = 8'h00;
	ram[7984] = 8'h00;	ram[7985] = 8'h00;	ram[7986] = 8'h00;	ram[7987] = 8'h00;
	ram[7988] = 8'h00;	ram[7989] = 8'h00;	ram[7990] = 8'h00;	ram[7991] = 8'h00;
	ram[7992] = 8'h00;	ram[7993] = 8'h00;	ram[7994] = 8'h00;	ram[7995] = 8'h00;
	ram[7996] = 8'h00;	ram[7997] = 8'h00;	ram[7998] = 8'h00;	ram[7999] = 8'h00;
	ram[8000] = 8'h00;	ram[8001] = 8'h00;	ram[8002] = 8'h00;	ram[8003] = 8'h00;
	ram[8004] = 8'h00;	ram[8005] = 8'h00;	ram[8006] = 8'h00;	ram[8007] = 8'h00;
	ram[8008] = 8'h00;	ram[8009] = 8'h00;	ram[8010] = 8'h00;	ram[8011] = 8'h00;
	ram[8012] = 8'h00;	ram[8013] = 8'h00;	ram[8014] = 8'h00;	ram[8015] = 8'h00;
	ram[8016] = 8'h00;	ram[8017] = 8'h00;	ram[8018] = 8'h00;	ram[8019] = 8'h00;
	ram[8020] = 8'h00;	ram[8021] = 8'h00;	ram[8022] = 8'h00;	ram[8023] = 8'h00;
	ram[8024] = 8'h00;	ram[8025] = 8'h00;	ram[8026] = 8'h00;	ram[8027] = 8'h00;
	ram[8028] = 8'h00;	ram[8029] = 8'h00;	ram[8030] = 8'h00;	ram[8031] = 8'h00;
	ram[8032] = 8'h00;	ram[8033] = 8'h00;	ram[8034] = 8'h00;	ram[8035] = 8'h00;
	ram[8036] = 8'h00;	ram[8037] = 8'h00;	ram[8038] = 8'h00;	ram[8039] = 8'h00;
	ram[8040] = 8'h00;	ram[8041] = 8'h00;	ram[8042] = 8'h00;	ram[8043] = 8'h00;
	ram[8044] = 8'h00;	ram[8045] = 8'h00;	ram[8046] = 8'h00;	ram[8047] = 8'h00;
	ram[8048] = 8'h00;	ram[8049] = 8'h00;	ram[8050] = 8'h00;	ram[8051] = 8'h00;
	ram[8052] = 8'h00;	ram[8053] = 8'h00;	ram[8054] = 8'h00;	ram[8055] = 8'h00;
	ram[8056] = 8'h00;	ram[8057] = 8'h00;	ram[8058] = 8'h00;	ram[8059] = 8'h00;
	ram[8060] = 8'h00;	ram[8061] = 8'h00;	ram[8062] = 8'h00;	ram[8063] = 8'h00;
	ram[8064] = 8'h00;	ram[8065] = 8'h00;	ram[8066] = 8'h00;	ram[8067] = 8'h00;
	ram[8068] = 8'h00;	ram[8069] = 8'h00;	ram[8070] = 8'h00;	ram[8071] = 8'h00;
	ram[8072] = 8'h00;	ram[8073] = 8'h00;	ram[8074] = 8'h00;	ram[8075] = 8'h00;
	ram[8076] = 8'h00;	ram[8077] = 8'h00;	ram[8078] = 8'h00;	ram[8079] = 8'h00;
	ram[8080] = 8'h00;	ram[8081] = 8'h00;	ram[8082] = 8'h00;	ram[8083] = 8'h00;
	ram[8084] = 8'h00;	ram[8085] = 8'h00;	ram[8086] = 8'h00;	ram[8087] = 8'h00;
	ram[8088] = 8'h00;	ram[8089] = 8'h00;	ram[8090] = 8'h00;	ram[8091] = 8'h00;
	ram[8092] = 8'h00;	ram[8093] = 8'h00;	ram[8094] = 8'h00;	ram[8095] = 8'h00;
	ram[8096] = 8'h00;	ram[8097] = 8'h00;	ram[8098] = 8'h00;	ram[8099] = 8'h00;
	ram[8100] = 8'h00;	ram[8101] = 8'h00;	ram[8102] = 8'h00;	ram[8103] = 8'h00;
	ram[8104] = 8'h00;	ram[8105] = 8'h00;	ram[8106] = 8'h00;	ram[8107] = 8'h00;
	ram[8108] = 8'h00;	ram[8109] = 8'h00;	ram[8110] = 8'h00;	ram[8111] = 8'h00;
	ram[8112] = 8'h00;	ram[8113] = 8'h00;	ram[8114] = 8'h00;	ram[8115] = 8'h00;
	ram[8116] = 8'h00;	ram[8117] = 8'h00;	ram[8118] = 8'h00;	ram[8119] = 8'h00;
	ram[8120] = 8'h00;	ram[8121] = 8'h00;	ram[8122] = 8'h00;	ram[8123] = 8'h00;
	ram[8124] = 8'h00;	ram[8125] = 8'h00;	ram[8126] = 8'h00;	ram[8127] = 8'h00;
	ram[8128] = 8'h00;	ram[8129] = 8'h00;	ram[8130] = 8'h00;	ram[8131] = 8'h00;
	ram[8132] = 8'h00;	ram[8133] = 8'h00;	ram[8134] = 8'h00;	ram[8135] = 8'h00;
	ram[8136] = 8'h00;	ram[8137] = 8'h00;	ram[8138] = 8'h00;	ram[8139] = 8'h00;
	ram[8140] = 8'h00;	ram[8141] = 8'h00;	ram[8142] = 8'h00;	ram[8143] = 8'h00;
	ram[8144] = 8'h00;	ram[8145] = 8'h00;	ram[8146] = 8'h00;	ram[8147] = 8'h00;
	ram[8148] = 8'h00;	ram[8149] = 8'h00;	ram[8150] = 8'h00;	ram[8151] = 8'h00;
	ram[8152] = 8'h00;	ram[8153] = 8'h00;	ram[8154] = 8'h00;	ram[8155] = 8'h00;
	ram[8156] = 8'h00;	ram[8157] = 8'h00;	ram[8158] = 8'h00;	ram[8159] = 8'h00;
	ram[8160] = 8'h00;	ram[8161] = 8'h00;	ram[8162] = 8'h00;	ram[8163] = 8'h00;
	ram[8164] = 8'h00;	ram[8165] = 8'h00;	ram[8166] = 8'h00;	ram[8167] = 8'h00;
	ram[8168] = 8'h00;	ram[8169] = 8'h00;	ram[8170] = 8'h00;	ram[8171] = 8'h00;
	ram[8172] = 8'h00;	ram[8173] = 8'h00;	ram[8174] = 8'h00;	ram[8175] = 8'h00;
	ram[8176] = 8'h00;	ram[8177] = 8'h00;	ram[8178] = 8'h00;	ram[8179] = 8'h00;
	ram[8180] = 8'h00;	ram[8181] = 8'h00;	ram[8182] = 8'h00;	ram[8183] = 8'h00;
	ram[8184] = 8'h00;	ram[8185] = 8'h00;	ram[8186] = 8'h00;	ram[8187] = 8'h00;
	ram[8188] = 8'h00;	ram[8189] = 8'h00;	ram[8190] = 8'h00;	ram[8191] = 8'h00;
end

//-----------------------------------------------------------------------------
always @(posedge clk)
begin
    if (we)
    begin
        ram[addr] <= din;
        dout <= din;
    end
    else
        dout <= ram[addr];
end

endmodule
//-----------------------------------------------------------------------------
