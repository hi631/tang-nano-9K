//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Fri Sep 30 16:21:12 2022

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire [29:0] prom_inst_4_dout_w;
wire [29:0] prom_inst_5_dout_w;
wire [29:0] prom_inst_6_dout_w;
wire [29:0] prom_inst_7_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h33333333333333333333333333333333B333333333333333333B3B3B3B3B3B33;
defparam prom_inst_0.INIT_RAM_01 = 256'h00000000000280888C84343C4140155340D055403CA14541FFDA7C0010434008;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h43350300C400CC4307D40C3004C31184343C334C310B032CD00C30000C80C000;
defparam prom_inst_0.INIT_RAM_05 = 256'hEB60D8B4CFC4F4D33AD4C0F3D31CEECCB903D834D4C0F3D31CC4F6D3434D0B0F;
defparam prom_inst_0.INIT_RAM_06 = 256'hB1B381B3831009321B400D6CC434601892208C888402C22402C22402C2004261;
defparam prom_inst_0.INIT_RAM_07 = 256'h0C08AB4C26B4020A263B080ED0C3B42D0B40000D10CC98ED0088089AD2F50D1B;
defparam prom_inst_0.INIT_RAM_08 = 256'h8918C00C4818E9B2CC03A393932C9A2283028022608A0C0A00898308302260C2;
defparam prom_inst_0.INIT_RAM_09 = 256'h020226B6302ED826E009AA08F00D000DA88C542C3000D8F80E380E0308EAE30C;
defparam prom_inst_0.INIT_RAM_0A = 256'h02263383C000CEC88C9AAA822AA634262D2248288AE1C910040810A00834AAA6;
defparam prom_inst_0.INIT_RAM_0B = 256'h088C00002AE280EB0A3030EDEA0088FB430E1C80800C02C88E980A0898202222;
defparam prom_inst_0.INIT_RAM_0C = 256'h00C0418843E0C8083C2B0B00203C010F20203C0103202041008F044EE1C0E00A;
defparam prom_inst_0.INIT_RAM_0D = 256'h0F0E30CC23A00401058CBB50C2C892482A0080F060015A4030282BED4ABA2A80;
defparam prom_inst_0.INIT_RAM_0E = 256'hDE1CE98A0B000B48AD0022C0822A8022BB500B70400A810C18FB60A90CC910CB;
defparam prom_inst_0.INIT_RAM_0F = 256'h102020BC0B8272000B070F08F08F00C308088882A3A62988AAAA0AA1BC400E00;
defparam prom_inst_0.INIT_RAM_10 = 256'h08A8E90B82820A90B82062020E0AA8288CBBB33BBBBB33BBBBBBBBB330C12321;
defparam prom_inst_0.INIT_RAM_11 = 256'h882028028C08B82286C0B0B030B22A8283022E82620082200AA402282A88802C;
defparam prom_inst_0.INIT_RAM_12 = 256'h8C8210400083C3008322288AAA008A338244B22E3C03200000008C8C00220E00;
defparam prom_inst_0.INIT_RAM_13 = 256'h228A280088C840A3030020088088B828F824FB60C083228C0BB5030730F00002;
defparam prom_inst_0.INIT_RAM_14 = 256'h2C0C8820830000082B038300C0BCC8B808A38C882E228088303000240E08C420;
defparam prom_inst_0.INIT_RAM_15 = 256'h202280220C8CC0938822008832C8C882080128BB60088B828CC8848B02200883;
defparam prom_inst_0.INIT_RAM_16 = 256'h220E0220200018AC8E0824801202ED4022282E022D8038B402AD8C0A2C38B302;
defparam prom_inst_0.INIT_RAM_17 = 256'hED0E002D0A8E000ADB4382888822228C88208E000208A8C1030098C20B8B4883;
defparam prom_inst_0.INIT_RAM_18 = 256'h02102AC2022420022A802AA20AD80238108E423B8002B782B621221020E00282;
defparam prom_inst_0.INIT_RAM_19 = 256'h2008300080088280230224A301028B0220E086084802088032C0B02F0E00AF03;
defparam prom_inst_0.INIT_RAM_1A = 256'h3B48B828C8890300022920823230020204012C0220012C01248088022800A089;
defparam prom_inst_0.INIT_RAM_1B = 256'h0E08F8A889A0281040220E0280822BC0E08080410020228C28E1C83002E0BB40;
defparam prom_inst_0.INIT_RAM_1C = 256'hC1D7036CF03C8D12060608880B08080802300836F0E08300AAA882AA02228ABC;
defparam prom_inst_0.INIT_RAM_1D = 256'h62188883604ECCCCCECEECECEED8B4968B4015B400D6CC43446E810022101028;
defparam prom_inst_0.INIT_RAM_1E = 256'h01888876088762188887608876018888B608876218888B608876018888360887;
defparam prom_inst_0.INIT_RAM_1F = 256'h08B400180621812F404B98880600000041D00874082D008B4080D00874008876;
defparam prom_inst_0.INIT_RAM_20 = 256'h80623180188F6874000D02834040018801000C60184223108420004040008C81;
defparam prom_inst_0.INIT_RAM_21 = 256'h2DB002DB001D8002D9180C10042200D88B420006218008F4006F0B0AE0210801;
defparam prom_inst_0.INIT_RAM_22 = 256'h001D00403D8004008F4000000010203D8080808040088B688840003D2002D900;
defparam prom_inst_0.INIT_RAM_23 = 256'h81D808080806080D8006080601D88F40010001D00403D8004080601D88F40010;
defparam prom_inst_0.INIT_RAM_24 = 256'h0042180600D8004082D8006081D8006081D8006081D80060080401D886080060;
defparam prom_inst_0.INIT_RAM_25 = 256'h00180C40001D00180C600D88362310188F6004018800C403D8018004003188B4;
defparam prom_inst_0.INIT_RAM_26 = 256'h320603D80188010042F01D80060800100403D8080808060042318834088C400D;
defparam prom_inst_0.INIT_RAM_27 = 256'h98880001000403D8834221342108400402C0802CC0108360041834C840318800;
defparam prom_inst_0.INIT_RAM_28 = 256'h04218880D008F40421000004002108B6B405053D7F4180000B42189888020318;
defparam prom_inst_0.INIT_RAM_29 = 256'h880100401D80D01001880108C4022004222231808818B6004000621888834018;
defparam prom_inst_0.INIT_RAM_2A = 256'h801800100400062101801806000680032060100040D88010042108018180602D;
defparam prom_inst_0.INIT_RAM_2B = 256'h2108760420062188B028B300601D8018880108C4220042222318081806000210;
defparam prom_inst_0.INIT_RAM_2C = 256'hD000603D08B6040043D80180600042108B4022004202231880603D8018801004;
defparam prom_inst_0.INIT_RAM_2D = 256'h008818F6B400D0274034C1800D600D03423108018080C62006088C6000600403;
defparam prom_inst_0.INIT_RAM_2E = 256'hCC8D0D433BF03198C2F16205014034F888C62000188888C60006042108042004;
defparam prom_inst_0.INIT_RAM_2F = 256'h1804018033BE3084C32D4B513C8000C8E478CCEE207471C71C72721288C476E5;
defparam prom_inst_0.INIT_RAM_30 = 256'h00CB4208B2D002CB40B01D131D800004008418B6C0BC80B881804118C4218C41;
defparam prom_inst_0.INIT_RAM_31 = 256'h48842CB42000203006030A30100CB4218802232D88400800CB42208800CB4208;
defparam prom_inst_0.INIT_RAM_32 = 256'h9D170785184810412103004818760684C2122D8880202D8040C202D884288042;
defparam prom_inst_0.INIT_RAM_33 = 256'h00000028000000002B32C170789682AAAAAAAAAAA40690AEAAAAAAAAAA046900;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h777777777777777777777777777777773777777777777777BBB3F73B7FB3F7FF;
defparam prom_inst_1.INIT_RAM_01 = 256'h000000000003038F0F8F37334201C40B0EC31175C30C3132DDC516DE28B31127;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'hBB39EB0CF683CF73E367FF3FFFFFFD8F3733F78F36C3FFCDE90C30D0CF0FF000;
defparam prom_inst_1.INIT_RAM_05 = 256'hCF81E4785FF6F9E3B0D8EBF7E36ECCCC834BE4B8D8EBF7E360D9F8EB83BEC3EF;
defparam prom_inst_1.INIT_RAM_06 = 256'hB1FF41BF03DCC2FF13840E4CD038742C55908F0F8F3DBECBAF75E71D3CC0C0F0;
defparam prom_inst_1.INIT_RAM_07 = 256'hCF2C6F87B7F83B6B17B42C5FE017FAFE3FAE6B2E7D075CFE02EE2C5CE104CE17;
defparam prom_inst_1.INIT_RAM_08 = 256'h70DED0C1B8EC75F100C0E04030B05DFFF33BC0BD77EFCCEF02F5C3EF3CB170FB;
defparam prom_inst_1.INIT_RAM_09 = 256'h0B8B17FAF8BFEB17F045FD0CF02E002ED940044F30001EF8010702002C66F1C3;
defparam prom_inst_1.INIT_RAM_0A = 256'h4F17B08005040E2FC45FFF4BBFD7B9FB3E77806FFCC1F0E3338840A31BBA3317;
defparam prom_inst_1.INIT_RAM_0B = 256'h6D845B50DFC3CF2F8F3E18CE7C034B3F8FC50F43588FC32FC65C3F2C5CB4BBFF;
defparam prom_inst_1.INIT_RAM_0C = 256'h14350DDB0CC3FC340E3F8FF0D3CC0903F0D3CE398BF0D079C3CFC433E3F5C00B;
defparam prom_inst_1.INIT_RAM_0D = 256'h4334004FB11CA50125EEFFBF30740E307B41CF3C304C0B4040EF74FEFCCABB1D;
defparam prom_inst_1.INIT_RAM_0E = 256'hEF3F35FFFF800FAEFE3F3FC2EF3FF0FD7FBC1FAE44050D4F5EFFBFF8C0F0CC3C;
defparam prom_inst_1.INIT_RAM_0F = 256'hD0FE32FF2FC33E032F07FFFEFFDFF8F530CDDDEFB1976FFFCFBBEE51FEB0C232;
defparam prom_inst_1.INIT_RAM_10 = 256'h2DB93CCF8B83D3CDFCB53131D393FC704F733FB733333F3333F33B33F180D1F0;
defparam prom_inst_1.INIT_RAM_11 = 256'hFF31F0CFCF0CF833CFE0FCFE3C3E0D474F0B74C3374C53740EF38F2C32CCFABE;
defparam prom_inst_1.INIT_RAM_12 = 256'hC3034C0E0ED3F3C7F3C333C57770FD3F4333433D14D03C033C30FFCF33FFCE1B;
defparam prom_inst_1.INIT_RAM_13 = 256'hFF4D1400CCF4F3E38BC3F03430FCF8F378337FBFCCD033020FFBC34BFC3C3C33;
defparam prom_inst_1.INIT_RAM_14 = 256'hF340CDBBE3C44703FCD303C3E3D538F00FCD80CD3BFF00CF3E304857CE1CF41C;
defparam prom_inst_1.INIT_RAM_15 = 256'h70FF4033CF03E3CD4CFF00CF3D340CDBEFC2F0FFBD2DFFCF3434C3FF33700CF3;
defparam prom_inst_1.INIT_RAM_16 = 256'hBB0C1F31FCC70017C1785F8C2F43FE34B7F03D033EFC3CF8D0FEBE3D1F7CF333;
defparam prom_inst_1.INIT_RAM_17 = 256'hFE3F003E3E3F003FEF8F4F0FCC77FF00CDBFCE1845B4F4F2F3C7E00FECCFBFD0;
defparam prom_inst_1.INIT_RAM_18 = 256'h4600F24F4FACF30FFCF013533FECCF1CC3C4FF7CF00FF8CFF830F37CF0F1E343;
defparam prom_inst_1.INIT_RAM_19 = 256'hB09F3851CC3FE4D1BF0B73373BE7073FBCF1539D7C773FD10FF3C0DFCE1DDFF3;
defparam prom_inst_1.INIT_RAM_1A = 256'h33BCF8F40CC033C7ABF8F80C3C3052174FC4E3C4E3C5E7C7E383EE3FBC32C5FC;
defparam prom_inst_1.INIT_RAM_1B = 256'hCE13FFEFE3ECFC4C0DFFCE1FB3EFBBFCD1F3F13038B6BB04F8C1F73073C0FF8F;
defparam prom_inst_1.INIT_RAM_1C = 256'hF3EF3785DE731CD9673A3EF607C604C40F3E1300FCF184F3BB2FFEEDCFF2CB3F;
defparam prom_inst_1.INIT_RAM_1D = 256'hB32C844FBC0DEEDCDFDCCDFDEDD8789407BE293840E4CD03845EE42C32836CEB;
defparam prom_inst_1.INIT_RAM_1E = 256'h1284007BC847B32C8447BCC8B8320C88FBC0C791240CCFBC40BA128400FBC847;
defparam prom_inst_1.INIT_RAM_1F = 256'h407A2200401252BDACAF240CC200130002E0007B013EC147B063EC28BB0040BA;
defparam prom_inst_1.INIT_RAM_20 = 256'h4811120C0447A0BB0D1EC343B00000C0804C0410280301080B112000103E8780;
defparam prom_inst_1.INIT_RAM_21 = 256'h3ED102EC213EC322EC000488423001E00F802AA2108040F9003DEFF3CF30C880;
defparam prom_inst_1.INIT_RAM_22 = 256'h211EC8333EC8810CCF8022022200012E40C848C80000C7B444B2112E0320ED03;
defparam prom_inst_1.INIT_RAM_23 = 256'hC2E008808883013E488208C202ECCF82204102E84223E88810C0311E00F92204;
defparam prom_inst_1.INIT_RAM_24 = 256'h8800044003E08800C3E08820C1E08820C0E08820C2E0882008C003E042808810;
defparam prom_inst_1.INIT_RAM_25 = 256'hC2008C32110E400004133EC8F8210E0CCFB003320C4C4221EC204001301000F8;
defparam prom_inst_1.INIT_RAM_26 = 256'h1E0003E820C0804013DF1EC8830008084220E800888082002110003B88C4112E;
defparam prom_inst_1.INIT_RAM_27 = 256'h4C347220433100E007B21079104C920033CF103C7400C3B00328788C23100CFA;
defparam prom_inst_1.INIT_RAM_28 = 256'h020083E3ECC83B011044B600321040F9FA0156C040818822038004C43882210C;
defparam prom_inst_1.INIT_RAM_29 = 256'h4880C8331EA0EC0C00C0804042030201202310C40A087B002320330C844FA000;
defparam prom_inst_1.INIT_RAM_2A = 256'h48000808430200304000044000018F11E0320E0000E048084330C8808088110E;
defparam prom_inst_1.INIT_RAM_2B = 256'h30C8F80102021084F3F4F1C0110E00004880C841012023130100860CC212E208;
defparam prom_inst_1.INIT_RAM_2C = 256'hE400111E403B010012E800C033201000CB8301202023010000332EE208C800C0;
defparam prom_inst_1.INIT_RAM_2D = 256'h3D3400397A07EA03A879C8801C230E0BA110C88048CC40220380441120308222;
defparam prom_inst_1.INIT_RAM_2E = 256'hCC5202C0008501018C40B310441101F0484222D8040C48422203021048C03002;
defparam prom_inst_1.INIT_RAM_2F = 256'hDCB63D03000B000111004011310444C100B0CC7743C471C71C71C3CC8B795406;
defparam prom_inst_1.INIT_RAM_30 = 256'h0443A208D0E202438830714DE10031C600031CFBFEF782F3810773D4B43D8352;
defparam prom_inst_1.INIT_RAM_31 = 256'h0088343B003F001C0A012912C0843B000423010E44B1808C438130480443A388;
defparam prom_inst_1.INIT_RAM_32 = 256'hDD3B90891E381002F003048C10FAC88A43283E8411132EC4100B02E00A30C0B3;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000002800000000380203B90AFCCFFFFFFFFFFF500D7BD2FFFFFFFFFF0CD40B;
defparam prom_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h777777777777777777777777777777773777777777777777B777333FFBBB773F;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000000000010B0343433733C3C3FFF8CE33FD70FFAD7FF34470C3FE3CF0D020;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_04 = 256'hD33FC70CFF03CFC1C33FFF7FFFF3FF03373347CF33C3FFCDFE0C30D0CFC7F000;
defparam prom_inst_2.INIT_RAM_05 = 256'h73E3F03CBDFFFDF700CDC8C7F330C8C83C0FF0FCCDC8C7F33CCDFCF3E7CFC3FF;
defparam prom_inst_2.INIT_RAM_06 = 256'h937D834D83FFC0CCB3CC0FCC703CD0087D4183C3C30C30D34D38E3CF3CC00F30;
defparam prom_inst_2.INIT_RAM_07 = 256'hC3086FCF2DFCF2421D580803F000FCFFBFCE232F4C0B763F04894877F1FCCF39;
defparam prom_inst_2.INIT_RAM_08 = 256'h34F543C1F7C8B75102C43464842074E3B332C92DDF9ECCCB24B743C83C21DC32;
defparam prom_inst_2.INIT_RAM_09 = 256'h42421DFFC423F31D7007780C4C2F002FD050001F0C0537725242509408B5D3C0;
defparam prom_inst_2.INIT_RAM_0A = 256'h521D5490005000088877AE122EDDBDEE0FEEC4BBBB12FCF313C0C0313FBFEEDD;
defparam prom_inst_2.INIT_RAM_0B = 256'h68003300C6118738C63E0C2F1903030FECC32F830B0FC60888770B0875292222;
defparam prom_inst_2.INIT_RAM_0C = 256'h08330EAFAC12F0300118CBD0C0C1188FD0C0C3080FD0C508C34FD07203F42042;
defparam prom_inst_2.INIT_RAM_0D = 256'h0330090F22D0201463768FCC227C8C3C0AC3830CA44C0A0023EBE03F318A2A8C;
defparam prom_inst_2.INIT_RAM_0E = 256'hF21F376E384103C8BFBB6E20823B802DCFDE0FDE01004C0F374FEC24D0FCCD08;
defparam prom_inst_2.INIT_RAM_0F = 256'hC12060BF48467D0348C7CFE8FE8FE0F43ACA8B82E29DB8BB92EECB735C72C0B2;
defparam prom_inst_2.INIT_RAM_10 = 256'h09E62CC8C28262CE842620342222ECA50F3773F3F777BB7777B77F7BB4C0C1C0;
defparam prom_inst_2.INIT_RAM_11 = 256'hAB102DD20119886612318C3D007E188A02026AA32A0D06A25AB35E386F99B221;
defparam prom_inst_2.INIT_RAM_12 = 256'h47068C0C0CA3F000B0F6A8906640893C4A33066028E03C834C32834F10EAC003;
defparam prom_inst_2.INIT_RAM_13 = 256'h2298411098F834908FC368347D9A806384A38FECCDA066C318FCD00BC03C343A;
defparam prom_inst_2.INIT_RAM_14 = 256'hE302AAAFA0C00303E0C043C3338A36842B8E02AA6A2250983E080823C304F20D;
defparam prom_inst_2.INIT_RAM_15 = 256'hA12204260F03038E992250983F382AAAF808E28FEE2AB80E3935808B36A90983;
defparam prom_inst_2.INIT_RAM_16 = 256'hAAC202202CC30007007403C08ECA3FB8AAEC60023FF438FED1BFF3382F78B336;
defparam prom_inst_2.INIT_RAM_17 = 256'h3FB3040F39310438FFEC4E4B592222C198A38208C038E0F4F04088526B83FBB0;
defparam prom_inst_2.INIT_RAM_18 = 256'h4300205242012B0EABA10E0E38F0CE04C381BE2BA10E3F8E3FE8FE0D2C300686;
defparam prom_inst_2.INIT_RAM_19 = 256'h201B0811BD0894B1A20263A730E6033E2C105299343648B00E0380CFC30C8FF0;
defparam prom_inst_2.INIT_RAM_1A = 256'h0BF984E4199030032229ACAC3E0010068384C7C4C705C744C3478A0E203485B8;
defparam prom_inst_2.INIT_RAM_1B = 256'hC107FBB8A4B9288C0CEAC202648E23FC10648230312222C12031F70C36118FEF;
defparam prom_inst_2.INIT_RAM_1C = 256'h30F333C8CC334CFF1D3308B503D200D1D23C2300FC3088EBEAF8AFA992E38EBF;
defparam prom_inst_2.INIT_RAM_1D = 256'hE01C4C4BEC0DCECCDFCCDFEEDDF83C3D47FD133CC0FCC703CCC480E3480F0CC3;
defparam prom_inst_2.INIT_RAM_1E = 256'h11C4C4FEC887D318080FEC447D318C4CFEC407C214C08FEC007F210808BECCC7;
defparam prom_inst_2.INIT_RAM_1F = 256'h403D03084101010FD043B08C4331100002FC14FC0A3F03CBC002F0147C00CC7E;
defparam prom_inst_2.INIT_RAM_20 = 256'h0C3101840083CCFC043F0247C03000C040C000031432200847311030022C8F00;
defparam prom_inst_2.INIT_RAM_21 = 256'h0F3110F3223F3332F3040040400033F003D0155010040CBF000FC3B4EE104C40;
defparam prom_inst_2.INIT_RAM_22 = 256'h001FC0312F80C308C7D21120230C231F0804404C300C83CC0471311FB221F303;
defparam prom_inst_2.INIT_RAM_23 = 256'h83F4844804C20B1F00C1040021F08BC030C111F04022FC0C3000311F08BF030C;
defparam prom_inst_2.INIT_RAM_24 = 256'h0C100C4320FC0C3042F40C10E2FC0C1042F40C10E1FC0C1000C313F800CC0C30;
defparam prom_inst_2.INIT_RAM_25 = 256'h43044002020F8300C0301F447D100404CBC8C12148440132F930000213004CFE;
defparam prom_inst_2.INIT_RAM_26 = 256'h3C0210FC308C408C20FC1F40C30C8408C202F488480CC0000300C47D4880133F;
defparam prom_inst_2.INIT_RAM_27 = 256'hCCB0BC30433331F043F30036104C610230CB710CF40083F000103DCC220048B3;
defparam prom_inst_2.INIT_RAM_28 = 256'h82000B10F0E83C0030C4310120200CBC7C02FABBBBAB871107D00C04F8013004;
defparam prom_inst_2.INIT_RAM_29 = 256'h0040C0313F23F00C0004400800322103230300000C087E0C001031008083F000;
defparam prom_inst_2.INIT_RAM_2A = 256'h0404040042310220C0800C4330C18BB3C0102E0022FCC408C030C4404008033F;
defparam prom_inst_2.INIT_RAM_2B = 256'h30407F021101204C32C033D0322F40000040C402211021233000CC0C4323F208;
defparam prom_inst_2.INIT_RAM_2C = 256'hF00C311F087C020010F0304402101304CFD210101102200C80102F0308840882;
defparam prom_inst_2.INIT_RAM_2D = 256'h2CF0043C3C46F02FC43CC4000C021F0BC300C44080840221010440021010C130;
defparam prom_inst_2.INIT_RAM_2E = 256'h88EE3A8EEEAF32AB8AA2A22B8AA22900000310C404C0CC0201018310C8410003;
defparam prom_inst_2.INIT_RAM_2F = 256'hFCBC2F4B33EA33CBFF2FCBB32E8CCC8FFBAC88AAA2BCA28A28A3B2ABB803ABBA;
defparam prom_inst_2.INIT_RAM_30 = 256'h0C03C14C00F41303DC3004000B8C22CF300B303CEC3F013B030BC2F4BE2F8BF2;
defparam prom_inst_2.INIT_RAM_31 = 256'h0844003F222C333D0510100114403E01CB20000F4C5284C803C318CC8403E144;
defparam prom_inst_2.INIT_RAM_32 = 256'hAA3AB98AAA80340110030400387C0504C8120F08C0121F80720811F4C5100460;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000000DAAAAAAAA2D1B43AB9380CEAAAAAAAAAAAFEAAABCAAAAAAAAAAFAABFA;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFF777777733333333F;
defparam prom_inst_3.INIT_RAM_01 = 256'h000000000003C0C4C4C433334040D5544D13554500000571001041033CF36214;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_04 = 256'hD339FC04D7C30D7103074F3DF4F3DD003333978C324BCF4CF60F3F008C87D000;
defparam prom_inst_3.INIT_RAM_05 = 256'hD3F1C83EDFC5FCF7D0C0F4F3F328CCCC14C7F07CCCF4F3F324CCFCC3134D4BDF;
defparam prom_inst_3.INIT_RAM_06 = 256'hC1F4D1C4D3581003132C0C4F303050805C004040408208208208208208000510;
defparam prom_inst_3.INIT_RAM_07 = 256'h8140778105781001153A4B45E235789E2783402E410F575E20840457E1540C9C;
defparam prom_inst_3.INIT_RAM_08 = 256'h4114C0600000F543A4611111010056EB3720D80D5BACDC8360357B4335015A10;
defparam prom_inst_3.INIT_RAM_09 = 256'h824015781405E01561C5710D502E942EDCE4B20D142154F01790140500F7F060;
defparam prom_inst_3.INIT_RAM_0A = 256'h011531E61804B7000C573D021DD5BBDE7EECD0F73673CC7400D4D0B531B9DDD5;
defparam prom_inst_3.INIT_RAM_0B = 256'h345B015084514111C5F36D6E16020117818A3C02034D41400D540B00541E2121;
defparam prom_inst_3.INIT_RAM_0C = 256'h18170731C552C02045314B008047098B00804709CB00854D41DF841342CD7015;
defparam prom_inst_3.INIT_RAM_0D = 256'h1720580C03D80615357F17805354D4146DDB0118D10ADCB53470E15E00471DD6;
defparam prom_inst_3.INIT_RAM_0E = 256'hE42C356DF5085F881E031D4012F3460D979A27934458054C57D7801044CC4449;
defparam prom_inst_3.INIT_RAM_0F = 256'h4421387A0501B306054B0F64F64F64DC197A7B83E395F4BB41CDC7754C406042;
defparam prom_inst_3.INIT_RAM_10 = 256'h01E61C79008E21C6540219112121CC994CFBBFF77BBB33BBBB7FBFBFBC6D6161;
defparam prom_inst_3.INIT_RAM_11 = 256'h6740210104245019004054B318F0294903C0C60309047E903EF128EEC3B3A114;
defparam prom_inst_3.INIT_RAM_12 = 256'h848887040463E140A12EEFA9A930BA354C006CE7242231C11007848D10D9D423;
defparam prom_inst_3.INIT_RAM_13 = 256'h21FA9630B8C840514F00EC1C4BBB94C054C05780CB02CE08257825CF10700C1E;
defparam prom_inst_3.INIT_RAM_14 = 256'h518B3BDF75084342C071C30043041F943B010B3BEE2130B8375C8C11D708D210;
defparam prom_inst_3.INIT_RAM_15 = 256'hC1218C2E0DC14301F82130B8341CB3BDF618CB97837B398C041FA4832EC30B83;
defparam prom_inst_3.INIT_RAM_16 = 256'hCED422022D000404404404018CCE5E0DECE4E6205E28B178B39E04383C70372E;
defparam prom_inst_3.INIT_RAM_17 = 256'h5E07017EB014217BC7810CC0FA2121CB38D3462D8110E4C075C08841FB9FBB12;
defparam prom_inst_3.INIT_RAM_18 = 256'h0004204142041B6CB7341E7E3BC0DEC0DB300E33341EF39EF0E44E401D7213C1;
defparam prom_inst_3.INIT_RAM_19 = 256'h2063502644484863D380C08F113D172C0D6061261C4908436C53080F870F4FB5;
defparam prom_inst_3.INIT_RAM_1A = 256'h5BB05CC8B3802143112408973658B609C4C844C8440844084443450D10206879;
defparam prom_inst_3.INIT_RAM_1B = 256'hD407FBB89010188704D9D502004D13ED6000421C1113DE041C73CB5C2E405783;
defparam prom_inst_3.INIT_RAM_1C = 256'h00F3332CCC330CDD0532047727472444013021D0F8600872FBB88BEC01EEECFE;
defparam prom_inst_3.INIT_RAM_1D = 256'hF3000CCBC12EEEEEDCCFFECCCFD0BC167BC50132C0C4F303074EE0001F800100;
defparam prom_inst_3.INIT_RAM_1E = 256'h3000CC7C58CFC3044007C1C0FD008440FC504FE10C884FC148FE200CC8BC548F;
defparam prom_inst_3.INIT_RAM_1F = 256'h0C7E0448C000000D00034840810110DD12F4447C113F044FC162F058BC1148FF;
defparam prom_inst_3.INIT_RAM_20 = 256'h8833000040CFCCBC902F140FCD0044C044480121080200488221110930100414;
defparam prom_inst_3.INIT_RAM_21 = 256'h2F1632F1631F1631F14CC144013200F4430111121080C43C5D0DC370DD20C444;
defparam prom_inst_3.INIT_RAM_22 = 256'h633FCC330FC110D4C3C040404042600F414141410DD04FC54833222F1522F162;
defparam prom_inst_3.INIT_RAM_23 = 256'h31FC1C1C1010571F01101C0103F403D0443413F84210F4110D48223FC83E0443;
defparam prom_inst_3.INIT_RAM_24 = 256'h5D230C4033FC110101F0110101F0110151F4110153F41101144222F81018110D;
defparam prom_inst_3.INIT_RAM_25 = 256'h1748C010033F174C81003FC0FD30404403D5D010C8801210F174C1110004C8BC;
defparam prom_inst_3.INIT_RAM_26 = 256'h105030F26488440C00DC3F01109CC4440110F414141411DD100488FC5441322F;
defparam prom_inst_3.INIT_RAM_27 = 256'h004440448DD230FC0310003F0040201120F4130F414C47D99108BC5D1104C040;
defparam prom_inst_3.INIT_RAM_28 = 256'h83104433F04CFC1330000112112080BCBC1155555541C30D17D208004487104C;
defparam prom_inst_3.INIT_RAM_29 = 256'h8844CC333F33F04374CC444C113131112123048C8044BD1D11112200CC87E048;
defparam prom_inst_3.INIT_RAM_2A = 256'h84488440C22110300437408111108421012310DD12F004484110844404C0021F;
defparam prom_inst_3.INIT_RAM_2B = 256'h000CFC12211030043D083D01103F77440044401020112322004CC0480301120C;
defparam prom_inst_3.INIT_RAM_2C = 256'hF811331F0C7C10DD22F074C0131112080FC220112232004880323F4444444C83;
defparam prom_inst_3.INIT_RAM_2D = 256'h10404CBCBC10F04BC130F4374F302F8BC304404449001201105441311105D320;
defparam prom_inst_3.INIT_RAM_2E = 256'h44551545555511554551511545511554001110044C88001211101200C4830DD0;
defparam prom_inst_3.INIT_RAM_2F = 256'h1005014011551145551545511544444555544455515451451451515555555555;
defparam prom_inst_3.INIT_RAM_30 = 256'h0403000880C03203003C55555580611601C45C30DC3714373500401004010040;
defparam prom_inst_3.INIT_RAM_31 = 256'h08C10132011301101130530504C031108402000C843004800333004CC4033008;
defparam prom_inst_3.INIT_RAM_32 = 256'h150015011450102C00BB201850BC404041010CC801212F88300722FC80008C00;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000000100000000011040015051040000000000500141140000000000001401;
defparam prom_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[29:0],dout[9:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 2;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h444444444444444444444444444444444444444444444444888888888888880C;
defparam prom_inst_4.INIT_RAM_01 = 256'h000000000000101010100303A0A2EAA8BA2EA9403CA14AB23B2DB6A31CF38000;
defparam prom_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_04 = 256'h0002D8080B400094200B130CF130CE9003030C83C004DC823443CC3000172000;
defparam prom_inst_4.INIT_RAM_05 = 256'h1844018403383220CC003830CC000C0D4280C544003830CC0B003030E00204C3;
defparam prom_inst_4.INIT_RAM_06 = 256'h4E404E404C242C00202C00833003A700A130C3C3C30C30C30C30C30C30F094B1;
defparam prom_inst_4.INIT_RAM_07 = 256'h700088B00A8B00002A0000822C0C88A2288FA2A2CA83A822C08380A822A800A4;
defparam prom_inst_4.INIT_RAM_08 = 256'h24A8000224883AA880008040C02CA9E7F700DA0EA79FDC03683A9801C002A600;
defparam prom_inst_4.INIT_RAM_09 = 256'h92532A88C932232A1D4AB27D0DE29DE2E020093E8DC028000088030008380002;
defparam prom_inst_4.INIT_RAM_0A = 256'hE02A082A08E201C800AB0EE20EEA88EC20ECDD3338073C7760DDDA77608AEEEA;
defparam prom_inst_4.INIT_RAM_0B = 256'h30D000B00E3720389CCF4D02F0C020088C1B73C00B70A28833A94B4CAA022220;
defparam prom_inst_4.INIT_RAM_0C = 256'hA00B07B1C6273C42037C9CF20803489CF00803489CF0038470DF02003732372C;
defparam prom_inst_4.INIT_RAM_0D = 256'h13004A122CE4220E1283088FB31CC60C8EDF2005CC001E073433C22234030EC4;
defparam prom_inst_4.INIT_RAM_0E = 256'h2073FA8E3858880822330E34C033840E0889688C80881AA0A8088F28032C0000;
defparam prom_inst_4.INIT_RAM_0F = 256'h0AA9D03C00DCCDC000DCCF70F70F770D1C7BBB896C6A383B00CEC78AA228012A;
defparam prom_inst_4.INIT_RAM_10 = 256'h4F6B047C933EB047893B0000B0F063ED30C44CC40444CC4444C8404488101814;
defparam prom_inst_4.INIT_RAM_11 = 256'h7377A8A8816305C8B00705CE058E30CEC353FBF90EC00EE835518C55C133B102;
defparam prom_inst_4.INIT_RAM_12 = 256'h224AC704041BE89E988EE3A2CC343B84DF330CE068CE02C1880BA2D1A0DCD363;
defparam prom_inst_4.INIT_RAM_13 = 256'hA838A03038022A30D8C2EC1223BB89F389F3888E4310CE79F888F4D8C1CC2C1E;
defparam prom_inst_4.INIT_RAM_14 = 256'h62033BDF741A1F40C8B058E317F82385F30E0338ECA8383A8741A1E2D07D1A8A;
defparam prom_inst_4.INIT_RAM_15 = 256'hC9A80E0EA12207CE3AA8383A862833BDF49EC3888F73381F3A2382A80CC383A8;
defparam prom_inst_4.INIT_RAM_16 = 256'hCED26AA6AD9D24A24A24A2C9EC8E223DCCECE168A225928897A2327963D2140C;
defparam prom_inst_4.INIT_RAM_17 = 256'h22337220B2206232088C9F323AAAA8033ADB616D5E24C308B45EA6083B083B10;
defparam prom_inst_4.INIT_RAM_18 = 256'h1E28AA088AA0835CF3340C1E320CDC0CDB822FF3340C830C81E89E8A8D069D5C;
defparam prom_inst_4.INIT_RAM_19 = 256'h2A734DF700AA3C23D353F3FFDCBD130C0D37B0FB122EAA334C17F0AFA37F6F34;
defparam prom_inst_4.INIT_RAM_1A = 256'h40BE09F433A0289F10AB08C6B349B67EA28C628C62CC62CC62C3430D0C002C30;
defparam prom_inst_4.INIT_RAM_1B = 256'hD17FF39ABC2080C704DCD17A820D0FCD17C2131C1321CE6089363345CE06088F;
defparam prom_inst_4.INIT_RAM_1C = 256'h281030000C0300E1CA2048BB0303000208C031DAFA070C40551A815608C554FC;
defparam prom_inst_4.INIT_RAM_1D = 256'h564995986821103321103111112D446A04418202C00833003A9128080D120892;
defparam prom_inst_4.INIT_RAM_1E = 256'h545515C6085C5545559C6089C5645559868C9C5645559868C9C5649559868C9C;
defparam prom_inst_4.INIT_RAM_1F = 256'h11C49184105414800520011110404602171805C60161A05860161A05868E85C4;
defparam prom_inst_4.INIT_RAM_20 = 256'h0D2748D98DD84D8600618018623E3801E8DD12344D13448D13747A3235405088;
defparam prom_inst_4.INIT_RAM_21 = 256'h71A3271A3271A3271A0C92C9D266771B000368E2749D9DC70600C0300C349DE8;
defparam prom_inst_4.INIT_RAM_22 = 256'h21711505713022045C5C1C1C1C8A12717070707228EC9C68C9155671A3271A32;
defparam prom_inst_4.INIT_RAM_23 = 256'h071F0F0F0B2200713022045057115C4C08821711505713022885057115C4C08A;
defparam prom_inst_4.INIT_RAM_24 = 256'h0E0349D3771B0228071F0228071F0220071F0220061F0228E413471E220F0228;
defparam prom_inst_4.INIT_RAM_25 = 256'h838C92266671A38C922771CDC6648889DC68E034999D22771A3828E004889D86;
defparam prom_inst_4.INIT_RAM_26 = 256'h422157183885E855140E617022485E859167170707072246324859C68C921671;
defparam prom_inst_4.INIT_RAM_27 = 256'h45050808200107145004540D141506205430054308815C60E205868E21481902;
defparam prom_inst_4.INIT_RAM_28 = 256'h52741036190D86E034D10BA37774D1C48660CD29BC221042E0504D45049B448D;
defparam prom_inst_4.INIT_RAM_29 = 256'hC9E8591661261D8808C9E899227267A2666648999C8DC646037A274D99DC6980;
defparam prom_inst_4.INIT_RAM_2A = 256'h5E885E855217A15498C085517460902426164202271C9E85932459E8D8592671;
defparam prom_inst_4.INIT_RAM_2B = 256'h4411866107A044150C050C260561808085E81522057A044454811C8150642141;
defparam prom_inst_4.INIT_RAM_2C = 256'h124603714DC7620202191801377A374D1853747A3777448DD1346180841E8D13;
defparam prom_inst_4.INIT_RAM_2D = 256'h400989C4C6031808620030808303610842489DE8A00D2277A200D2277A202277;
defparam prom_inst_4.INIT_RAM_2E = 256'h654850D4400EA320AC2C110050112134C921642E8555C92167A321645C916023;
defparam prom_inst_4.INIT_RAM_2F = 256'h2509425018C109084712D4BB03FA98B1448C8844E5059259E5970D1311400372;
defparam prom_inst_4.INIT_RAM_30 = 256'hDD20360448081120220DCE0502100408401021000C0380038A50942509425094;
defparam prom_inst_4.INIT_RAM_31 = 256'h00926200274027422264924989920274981274809D26049D202660499D202604;
defparam prom_inst_4.INIT_RAM_32 = 256'hAE09E0A004CC292024802E852904909202480055831641591601641592600926;
defparam prom_inst_4.INIT_RAM_33 = 256'h0000000C000000008C92209E0ECCAAAAAAAAAAA994620150AAAAAAAAA9122511;
defparam prom_inst_4.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[29:0],dout[11:10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 2;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h444444444444444444444444444444444444444444444444444444444444444C;
defparam prom_inst_5.INIT_RAM_01 = 256'h000000000000404040400000C0C03FFCD735FD4500000FC3733CF1CC00C0C000;
defparam prom_inst_5.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_04 = 256'hB44FC0000F0010C0142F104C3104C30000002CD3C2040CD10010C01000033000;
defparam prom_inst_5.INIT_RAM_05 = 256'hC4010040903D3D1405090D04EC2D01039AC4F041090D04EC2F093D34F4130413;
defparam prom_inst_5.INIT_RAM_06 = 256'h0F000F002C303C00300480C01203F380F013C3C3C30C30C30C30C30C30D0B1B0;
defparam prom_inst_5.INIT_RAM_07 = 256'h3080C4F00F4F00C33F3002053E014CD334CD9153442BFC53E00180FD33FC0030;
defparam prom_inst_5.INIT_RAM_08 = 256'h1C7CC8231C46BFD40020CCCC4C1CFCF3FF00F00FF3CFFC03C03FCC00C003F300;
defparam prom_inst_5.INIT_RAM_09 = 256'hC3C33F4CEC35333F0C0FF33F1CD3ECD3F002221E9CE03CCCC004C13087BC8823;
defparam prom_inst_5.INIT_RAM_0A = 256'h603F3000006128C4A8FF0C600CFF4CCC00CCFCF330B03CFF10FCF03F104DECFF;
defparam prom_inst_5.INIT_RAM_0B = 256'hF0F232100CA39030CE0FCF33F8401014CECE03400FF01208FBFF0E0CFC000000;
defparam prom_inst_5.INIT_RAM_0C = 256'h63230F33CCA03401063E80D0040A0C80D1040A0C80D2000010FF0100A030630C;
defparam prom_inst_5.INIT_RAM_0D = 256'h030000013EFC330003CF14CDB33CCD2C0CF3100CEC009C253C31C0533C0F3CCC;
defparam prom_inst_5.INIT_RAM_0E = 256'h3A03FFCC318C0000133F3CA0F0B30E0F14CE34CC200048033CD4CD2403140000;
defparam prom_inst_5.INIT_RAM_0F = 256'h02CFC03C008E0C400240CF30F30F3F0C3CF3332CCEFF303330CCCFC3D1142315;
defparam prom_inst_5.INIT_RAM_10 = 256'h0DE73CF2431E73CF243730807373C1EF33000808C0004800008408008E180C0C;
defparam prom_inst_5.INIT_RAM_11 = 256'h33D3C4ACC23B88EE73A3A40F240F30CCC383F3F73C400CC4F3334C31CF333309;
defparam prom_inst_5.INIT_RAM_12 = 256'h12CCCF0C4037D64F348CC304DCF0F30C8F33CCC301C60DC3493712C370CCF933;
defparam prom_inst_5.INIT_RAM_13 = 256'hCC3103F0F03D2B3200C1CC3D233308F308F314CD033CCCDB794CFE80E40C1C3C;
defparam prom_inst_5.INIT_RAM_14 = 256'hD33333FFFE4D4FC0C4E080C323F33308F30CF330CCCCF0F30FE4D4D3F93C3C4A;
defparam prom_inst_5.INIT_RAM_15 = 256'hCFCC3C3CC31323CC30CCF0F30D3B333FFCF0C314CFF3308F313303300CCF0F30;
defparam prom_inst_5.INIT_RAM_16 = 256'hCCF83C43CF0F3CD2CD2CD2CF0CCC533FCCCCC43C1330F04CC3D3383C03733C0C;
defparam prom_inst_5.INIT_RAM_17 = 256'h533730003134303004CE0F9230CCCCB333FFD83F0D38C334FE0F313C3300332C;
defparam prom_inst_5.INIT_RAM_18 = 256'h0F3CCD3CCCD3C3DC733C0C3EF00CFC8CF3212C733C0C030C03E4FE4ACF83FC0E;
defparam prom_inst_5.INIT_RAM_19 = 256'h0073ECFF00330CD3F303F3FFF4BF030C3FB3733B312CB313CC13F05F5B3FDF3E;
defparam prom_inst_5.INIT_RAM_1A = 256'hCCFFACF7331C16CF30C73CCF73ECFF3CD2CCD2CCD2CCD2CCD2C3030C04001CF0;
defparam prom_inst_5.INIT_RAM_1B = 256'hFB37FF331CD3C4CF0CCCFB3C4F0C07CFB34F133C3000CC53CCA033ECCCB394CF;
defparam prom_inst_5.INIT_RAM_1C = 256'h00300048000000304F10043C030000013CCD33F5F5B34CC0CC3303313CC31C7C;
defparam prom_inst_5.INIT_RAM_1D = 256'h030000CC1333332222221000033CC0FF5C430300480C01203DCC0434CCB00030;
defparam prom_inst_5.INIT_RAM_1E = 256'h30000CC13CCC030000CC13CCC030000CC1BCCC030000CC1BCCC030000CC13CCC;
defparam prom_inst_5.INIT_RAM_1F = 256'h0CC04C0C00303040CC103000002001303305CCC133306CCC1F3304CCC17CCCC0;
defparam prom_inst_5.INIT_RAM_20 = 256'hCC3200C40C8C08C133304CCC1017F0C0F0CC00330C33000CC3303C103300C040;
defparam prom_inst_5.INIT_RAM_21 = 256'h307E2307E2307E2307C8C0CCC33323053033244330CCC8C1300000000330CCF0;
defparam prom_inst_5.INIT_RAM_22 = 256'hE230CC32305301708C14D4D4D407C230535353501FC88C1F883332307E2307E2;
defparam prom_inst_5.INIT_RAM_23 = 256'h230131313101B2305301B8C3230C8C14C04E230CC3230530178C3230C8C14C04;
defparam prom_inst_5.INIT_RAM_24 = 256'hBC2208821301301B23013017230130132301301723013013C8C223010131301B;
defparam prom_inst_5.INIT_RAM_25 = 256'h6F04402221307F0480213044C22004084C1FC2108888021307F01FC2204084C1;
defparam prom_inst_5.INIT_RAM_26 = 256'h01021306F048F0882001301301348F088213013131310130120084C1F4802130;
defparam prom_inst_5.INIT_RAM_27 = 256'h040404C01001130440222001208421421000210004084C1B8104C1FC12008401;
defparam prom_inst_5.INIT_RAM_28 = 256'h813040030400C1C1104407C1111044C0C1037715C3974103C812040404812004;
defparam prom_inst_5.INIT_RAM_29 = 256'h04F0441030030404C004F044010113C1111100444400C130113C1004440C3404;
defparam prom_inst_5.INIT_RAM_2A = 256'h4F004F044013C110404C0441130000001010013003004F04401044F040441030;
defparam prom_inst_5.INIT_RAM_2B = 256'h1040C10013C110400000001010304C0C04F04400113C11111004440441000104;
defparam prom_inst_5.INIT_RAM_2C = 256'h01303330CCC101303304C004003C00000C00013C000010000400304C004F0040;
defparam prom_inst_5.INIT_RAM_2D = 256'h00040CC0C13304CC10000C4C003330CC000000F093000003C13000003C130033;
defparam prom_inst_5.INIT_RAM_2E = 256'h4585F00CCC8004000080449124444108C000301F0000C00003C100000C001303;
defparam prom_inst_5.INIT_RAM_2F = 256'h3C0F03C0100D54400090240010001231440DCE44353C71F71C773A10307220B0;
defparam prom_inst_5.INIT_RAM_30 = 256'hCC0031300004C0001001C041C3C0B02F02C0BC0000004C0043C0F03C0F03C0F0;
defparam prom_inst_5.INIT_RAM_31 = 256'h3083100032003201833023028CC00320C4C33000C83130CC0033130CCC003130;
defparam prom_inst_5.INIT_RAM_32 = 256'h100EC4AAD9CC38082028062CB80080813204C0CC4F3200C83133200C83130831;
defparam prom_inst_5.INIT_RAM_33 = 256'h0000000000000000C09020EC49CCAFFFFFFFFFFE4CB18C43FFFFFFFFFE23132C;
defparam prom_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[29:0],dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 2;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h000000000000000000000000000000000000000000000000000000000000000C;
defparam prom_inst_6.INIT_RAM_01 = 256'h0000000000022121212141410301C00200880160BEA96002D74515DC000208AA;
defparam prom_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_04 = 256'h2800DB082342E2086803028CB028C821414190220000ACA038A30CE0C22B2000;
defparam prom_inst_6.INIT_RAM_05 = 256'h200A320023323008AA022228C0060A0CB8E8C202022228C00002323888A200A3;
defparam prom_inst_6.INIT_RAM_06 = 256'hB883AC83AC0858C2C4481111E0470B040A60E3E3E38E38E38E38E38E38E83938;
defparam prom_inst_6.INIT_RAM_07 = 256'hB08C203130031380000984740C6500C0300E23408C130240C44A08000000110B;
defparam prom_inst_6.INIT_RAM_08 = 256'h38C03C4638C5302E58468282822802FBFF02FB2C0BEFFC0BECB02C0EC2300B03;
defparam prom_inst_6.INIT_RAM_09 = 256'hE2E20000DE2403006E803FBF5EC0EEC0CA9A4EAFDEC680382A682A0AC932EC46;
defparam prom_inst_6.INIT_RAM_0A = 256'h82000299A68A46889003ED812CC002DDB1DEDEBFF27B2CF7A3DEEFBFA302CCC0;
defparam prom_inst_6.INIT_RAM_0B = 256'hBFE4E3222C7B31F1ECCBDE50B080B1D00DEBB2808B82200893038B8800291212;
defparam prom_inst_6.INIT_RAM_0C = 256'h82330B31C47B280B77BDECA02C778AECA02C778AECA0228228FF2B1E7B297B4E;
defparam prom_inst_6.INIT_RAM_0D = 256'h3B08EB8224CE2B8A0803900E3B1EC63E6DEBB1DECA052F4AF47EC84038FB0CC4;
defparam prom_inst_6.INIT_RAM_0E = 256'h07B2B02DB5ED2C44803B0C78A33F0A2C900FB00E75268C0200100E083828C38E;
defparam prom_inst_6.INIT_RAM_0F = 256'hD1DEC8BC89ECC88089EC8FB8FB8FB82C2CF3332CC4C0B477A3FCCB202E344634;
defparam prom_inst_6.INIT_RAM_10 = 256'h8ACB0C75E22CB0C71E2B0E0EB0B0C2CF82444444444444444444444440A048C8;
defparam prom_inst_6.INIT_RAM_11 = 256'hBBBAD8DEE7B31ECCB07B1ECB9ECBBEECE0E2E3FB0C83ADC83731BE72EBFB3227;
defparam prom_inst_6.INIT_RAM_12 = 256'h23ECCF0808BBF9EB78EDDB76DEB03309EE33BEC780C80BC28C2F23C2F8EEE7A3;
defparam prom_inst_6.INIT_RAM_13 = 256'hDEB5EBB8302E37B9EC92CD2E3B775EE31EE3100E03BBECE3B100FDEC9EC92D2C;
defparam prom_inst_6.INIT_RAM_14 = 256'hA32FB3EFB9EAEB81E8F9E0827BB23B5EB78CEFB2DDDEB0330B9EAEA3E7AC2C8D;
defparam prom_inst_6.INIT_RAM_15 = 256'hEDDE2C0CC2237B8CB4DEB0330A3EFB3EFAEBEB500FB7B5EE323B5B780DEB0330;
defparam prom_inst_6.INIT_RAM_16 = 256'hECE7ADBADEEBBEE3EE3EE3EEBEED403EDEDED7BD003EF400FBC037BBB2BF740D;
defparam prom_inst_6.INIT_RAM_17 = 256'h4036B4B17A37B4B7200DEEE3B5DEDEEFB3EFA7AEEA3EF828F9EB720EB76C77BB;
defparam prom_inst_6.INIT_RAM_18 = 256'hEBBEDE0EEDE0EB9EBFFBEFACB72EED3EE78E3DBF79EDCB6DCAC8EC8DEE7AECEC;
defparam prom_inst_6.INIT_RAM_19 = 256'h1FBF9ABF4537AC3BE0E2E3FFE8FE3B0E2E6AB0B3323C77BB9E7BA0AFE6AFAFF9;
defparam prom_inst_6.INIT_RAM_1A = 256'h943B1AEEFB3839AB22DB0ECFBFDABAACE3ECE3ECE3ECE3ECE3E38B8E2A08AC3A;
defparam prom_inst_6.INIT_RAM_1B = 256'hE6ABF3336C20EECF08EEE6AD838E2BFE6A83BB3C2220ECE0EA6B2B9AAD6B100F;
defparam prom_inst_6.INIT_RAM_1C = 256'h070C1CE30EC3B0CA901888B3B93BBA3A0E0BB3EEFE6AECE1DCB747720EE72EBF;
defparam prom_inst_6.INIT_RAM_1D = 256'h1BB666E820E2222222222222210E40009402F84481111E04710298082D908423;
defparam prom_inst_6.INIT_RAM_1E = 256'hBB666E820EE81BB666E820EE81BB666E820EE81BB666E820EE81BB666E820EE8;
defparam prom_inst_6.INIT_RAM_1F = 256'h6E80803E6DBABBB02EEC06666D899A00FA082E820BA082E820BA082E8200EE81;
defparam prom_inst_6.INIT_RAM_20 = 256'hE2CB832832E82E820BA082E820C803E6832260CBB2F89832EC89A0E0CB86E183;
defparam prom_inst_6.INIT_RAM_21 = 256'hA083BA083BA083BA083E20B22C88BA020C78AAAC8B222E8200F06C1B078B2283;
defparam prom_inst_6.INIT_RAM_22 = 256'h3BA022CBA0200E02E808080808380BA020202020E00EE820EEC88BA083BA083B;
defparam prom_inst_6.INIT_RAM_23 = 256'hBA020202020E0BA0200E0E2CBA02E8080383BA022CBA0200E0E2CBA02E808038;
defparam prom_inst_6.INIT_RAM_24 = 256'h0CF8B22CBA0200E0BA0200E0BA0200E0BA0200E0BA0200E00E2CBA020E0200E0;
defparam prom_inst_6.INIT_RAM_25 = 256'h833EE0488BA0833E20CBA0EE80883832E820CFBB22220CBA0833200FB8032E82;
defparam prom_inst_6.INIT_RAM_26 = 256'h860CBA0833E28322CB07A0200E0E28322CBA020202020E0CF8832E820E20CBA0;
defparam prom_inst_6.INIT_RAM_27 = 256'hBE1E1803230FBA0EECC88BCF8B2ECA0CBB118BB11832E820CFBE820CF8832E1B;
defparam prom_inst_6.INIT_RAM_28 = 256'h2CBBE1BA08EE820F8B2E1A0C888B2E82820EAAFEAAACE7960838B2BE1E208832;
defparam prom_inst_6.INIT_RAM_29 = 256'hE28322CBA0BA083803E283220CB88A0C88888322283E8200F8A0CB9222E8383E;
defparam prom_inst_6.INIT_RAM_2A = 256'h283E28322F8A0C8B8380322CA00EE1B860CB8600FA0E28322F8B22838322CBA0;
defparam prom_inst_6.INIT_RAM_2B = 256'h8B2E820F8A0C8B2EC46EC460CBA0803EE283220F88A0C888883228322CB878B2;
defparam prom_inst_6.INIT_RAM_2C = 256'h0200FAA0EA820E00FA0803E2C8A0C8B2E83888A0C888883222CBA0803E28322C;
defparam prom_inst_6.INIT_RAM_2D = 256'h86183A82820A082820CF3B8033FAA0E838832283E0E20C8A0E0E20C8A0E00CAA;
defparam prom_inst_6.INIT_RAM_2E = 256'hBB8EA3A8888EEF33B8ACAAE2A8AAA14EA20CA8683222A20C8A0E0C8B2A2CA00E;
defparam prom_inst_6.INIT_RAM_2F = 256'h4A1284A1FC8BFEFC8BF2ECBBF2FFEFE288CBBB88AF2BEFAEBAEA2A23200332A3;
defparam prom_inst_6.INIT_RAM_30 = 256'hEE0C7A0283180A0C60C425200CA0284280A10AC706C182C180A1284A1284A128;
defparam prom_inst_6.INIT_RAM_31 = 256'h02AFA0C4BA84BA860FB82B82BEE0C7ABE80BB831EAFA02EE0C7BA02EEE0C7A02;
defparam prom_inst_6.INIT_RAM_32 = 256'hFBA1FC0CB28C0A93AA40088E0AC2AAAE0AB831EE83BAB0EAFA0BAB0EAFA02ABA;
defparam prom_inst_6.INIT_RAM_33 = 256'h00000000AAAAAAAA86D18A1FC3800AAAAAAAAAAABBFAFAA3AAAAAAAAAAFFAEFA;
defparam prom_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[29:0],dout[15:14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 2;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h4444444444444444444444444444444444444444444444444444444444444440;
defparam prom_inst_7.INIT_RAM_01 = 256'h0000000000011010101000004040155445115545000005400010410010404455;
defparam prom_inst_7.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_04 = 256'h5041D101074040441007100C3100C11000005440000410010440001090140000;
defparam prom_inst_7.INIT_RAM_05 = 256'h5444014640043510040004005004000010D0D144000400500400140010000403;
defparam prom_inst_7.INIT_RAM_06 = 256'h414C714C70D4D48D50140040100054405510D0D0D04104104104104104000534;
defparam prom_inst_7.INIT_RAM_07 = 256'h43C054430544304015140D45111544110441521149475551104140551154C054;
defparam prom_inst_7.INIT_RAM_08 = 256'h249440912480754540904040400055C73330CD0D571CCCC3343550C10F015430;
defparam prom_inst_7.INIT_RAM_09 = 256'hD0D015441D051015D345734CDD113D11D450D31E1D1014540144010040755091;
defparam prom_inst_7.INIT_RAM_0A = 256'h501514410450D50004571D510DD545DC13DCCD7B35750C3352CDC1735245DDD5;
defparam prom_inst_7.INIT_RAM_0B = 256'h78CD1250CD774335DD432C513447031441D3504B030011400757434055041010;
defparam prom_inst_7.INIT_RAM_0C = 256'h51270370C17504304771D410C0C740D410C0C740D410C00413CFC0317505741C;
defparam prom_inst_7.INIT_RAM_0D = 256'h03300D0001DD034011471441770DC12D5DCF031DD00F7CDF30F1F15104870DC0;
defparam prom_inst_7.INIT_RAM_0E = 256'h1750355D75D044C411070D741273430D544344414C44494054544114C0048C00;
defparam prom_inst_7.INIT_RAM_0F = 256'h84DCD03F01DD404301D40F30F30F300ECC37774DD1D5743712CDC35545209121;
defparam prom_inst_7.INIT_RAM_10 = 256'h41D70C35D01D70C35D0700207070D1DC00444444444444444444444444348484;
defparam prom_inst_7.INIT_RAM_11 = 256'h3334D48CD7775DDD70775D435D4370DDD1D0C7370D6C1DD43F706CF7C7B37007;
defparam prom_inst_7.INIT_RAM_12 = 256'h12DDC3000037E1D3749DD744DC703701DC006CD7540501E0480752C074CCC743;
defparam prom_inst_7.INIT_RAM_13 = 256'hDC750370350D2335D420DE0D27775DC05DC054410F36CDD7754431D41D420E0D;
defparam prom_inst_7.INIT_RAM_14 = 256'h121B37CF31D0D303C4B5D0007705275D3F01DB35DCDC7037031D0D12C74C0448;
defparam prom_inst_7.INIT_RAM_15 = 256'hCCDC1C0DC012770175DC7037012DB37CF1CDC754433F35DC052743703FC70370;
defparam prom_inst_7.INIT_RAM_16 = 256'hCDC74D34DCD35D52D52D52DCDCDD510CFCDDD74C510D314437110773507B303F;
defparam prom_inst_7.INIT_RAM_17 = 256'h510741137127413D0441DCD274DCDCDB37CF074CD12DC004B1D3510C7704F736;
defparam prom_inst_7.INIT_RAM_18 = 256'hD35DD50CDD50C71C7B304C1D3D0DCF4DCB112D7B304F430F41D49D48CC74CDDD;
defparam prom_inst_7.INIT_RAM_19 = 256'h31F31D33C8771C37C1D0C0CFC4BC033C0C747077012D37373C77001F874F1FB1;
defparam prom_inst_7.INIT_RAM_1A = 256'h14735DCDB35421D300D70DC37B1D334DD2DC12DC12DC12DC12D3034C04301C30;
defparam prom_inst_7.INIT_RAM_1B = 256'hC747F3775C10CDC300CCC74D430C07EC7443370C0001CDD0CD75071D1D775443;
defparam prom_inst_7.INIT_RAM_1C = 256'h30100014010040154500403743C340810C0370C5F874DC10FD7743F50CCF7C7E;
defparam prom_inst_7.INIT_RAM_1D = 256'h474111D45011111111111111111D4415344F010140040100045554040DC24892;
defparam prom_inst_7.INIT_RAM_1E = 256'h74111D450DD4474111D450DD4474111D450DD4474111D450DD4474111D450DD4;
defparam prom_inst_7.INIT_RAM_1F = 256'h1D44400D107474401D1001111044450035141D45075141D45075141D4500DD44;
defparam prom_inst_7.INIT_RAM_20 = 256'hD107401401D45D45075141D4500400D1C011100741344401D04470100741D040;
defparam prom_inst_7.INIT_RAM_21 = 256'h5153751537515375150D10C11044751100347FF044111D4500001004034411C0;
defparam prom_inst_7.INIT_RAM_22 = 256'h3751110751100101D44404040404075110101010100DD454DD04475153751537;
defparam prom_inst_7.INIT_RAM_23 = 256'h751101010101075110010D107511D444004375111075110010D107511D444004;
defparam prom_inst_7.INIT_RAM_24 = 256'h4C34411075110010751100107511001075110010751100100D10751101010010;
defparam prom_inst_7.INIT_RAM_25 = 256'h530DD0044751530D100751DD44440401D454C374111100751530100374001D45;
defparam prom_inst_7.INIT_RAM_26 = 256'h4100751530D1C01104035110014D1C01107511010101014C34401D454D100751;
defparam prom_inst_7.INIT_RAM_27 = 256'h4D0D04001233751DD0044403441D0500740047400401D454C34D454C34401D07;
defparam prom_inst_7.INIT_RAM_28 = 256'h1074D075149D4503441D070044441D45450155555555D34F0474414D0D144401;
defparam prom_inst_7.INIT_RAM_29 = 256'hD1C011075175140400D1C0110074470044444011140D45003470074111D4740D;
defparam prom_inst_7.INIT_RAM_2A = 256'h1C0D1C0113470044404001105001D07410074100351D1C01134411C040110751;
defparam prom_inst_7.INIT_RAM_2B = 256'h441D45034700441D001D00100751400DD1C01103447004444401140110743441;
defparam prom_inst_7.INIT_RAM_2C = 256'h11003751DD450100351400D104700441D474447004444401110751400D1C0110;
defparam prom_inst_7.INIT_RAM_2D = 256'h41040D454505141450000C40003751D4744011C0D0D10047010D100470100075;
defparam prom_inst_7.INIT_RAM_2E = 256'h5545515444455511545455515455515DD100741C0111D100470100441D105003;
defparam prom_inst_7.INIT_RAM_2F = 256'h1D0741D054455554455154555155555144455544551555555555151111511151;
defparam prom_inst_7.INIT_RAM_30 = 256'hDD003501400405001001454545D0741741D05D000100410041D0741D0741D074;
defparam prom_inst_7.INIT_RAM_31 = 256'h01D3500077407741037437434DD00374D4077400DD3501DD0037501DDD003501;
defparam prom_inst_7.INIT_RAM_32 = 256'h5505140555401D3474D4051D5D45D1D1074400DD437751DD3507751DD3501D35;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000400000000041100514444000000000000400105510000000000001005;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_pROM
