//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Mon Mar 14 11:49:20 2022

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h19E8ECAD26B498F0827FB7F37DC255DC05442097F095F0D02083000F000B000F;
defparam prom_inst_0.INIT_RAM_01 = 256'h85E91495614490480623426C240623422C355F42657D08ACDACF815BAD9D080A;
defparam prom_inst_0.INIT_RAM_02 = 256'h8A2137BA2895638219905E1990577D5DDDD608E15EB64F393E7896E4AB857A90;
defparam prom_inst_0.INIT_RAM_03 = 256'h75595EBBEEE1D57155C55793D947AF673923D9466767676494751454E8A27FFE;
defparam prom_inst_0.INIT_RAM_04 = 256'h8609D56C2F18CA7A4280808A4A86128138A1822256926A73391C93730FA5A9B8;
defparam prom_inst_0.INIT_RAM_05 = 256'h10001C0730F840000967C3CDD8784E2CE994972C60A1E0F87355871F38272272;
defparam prom_inst_0.INIT_RAM_06 = 256'h34C174F3D809BA45FD327672C0F926A8F098402AB92F6118111241C12AAAA5AA;
defparam prom_inst_0.INIT_RAM_07 = 256'h6FCB04FF8BF8E4E5DBC4D24959A8497E7F81E97F41C2CC14FDC9441F253EF119;
defparam prom_inst_0.INIT_RAM_08 = 256'h60D4700D93E6E098DD8082568D18FC96490754935E3D55F5A15A5EE72861F22E;
defparam prom_inst_0.INIT_RAM_09 = 256'hF6CDA66CF10594125101AE26A23262E8216FE2D908DC33F8E298306D5092FED4;
defparam prom_inst_0.INIT_RAM_0A = 256'h133A40CEB093667C7394CD0BC981D87B1B407CF6496F7C7C905C1AC7335A91A7;
defparam prom_inst_0.INIT_RAM_0B = 256'h68697EBE0140D824260423F4623909CD4D48649FF07C2A7F096ADE49BC6B26E7;
defparam prom_inst_0.INIT_RAM_0C = 256'hCF3E8366CF3D04C385EF8FAE9A707708C71055182674C8B85AECD14FC563C630;
defparam prom_inst_0.INIT_RAM_0D = 256'h5EE1B904D6827C242E91BA430C35C00000D4CF8B844E95CD8D885A404B232324;
defparam prom_inst_0.INIT_RAM_0E = 256'h89965C65997BB6D189269A69249A496CC85F63B49949A7BF2A17799D1161FEF8;
defparam prom_inst_0.INIT_RAM_0F = 256'h715768E5693687E9AF27597605F14B5C970505C931C954BD265B46DB41328794;
defparam prom_inst_0.INIT_RAM_10 = 256'h5696926B1DE79ADA6BFF683CCFB921EEF3B91A0EFC2EFFCAEEF04EFF95EFF4DA;
defparam prom_inst_0.INIT_RAM_11 = 256'h293A0ABEF82E09AE514152238A4AB92B69ED2AD229566B2E52979695A792FD67;
defparam prom_inst_0.INIT_RAM_12 = 256'h5D6E592DA5594822C26EE45FCB487BB189A599AA3B57740D69E49AFC5E234BB7;
defparam prom_inst_0.INIT_RAM_13 = 256'h4962E61A26D5255C4956A9224B92279AE63839EE42E527B092EED0B65578656A;
defparam prom_inst_0.INIT_RAM_14 = 256'hEE85F6DF93B9A5050171B18EE95D55E201987B2A6255EC673CBEE748ACA56E53;
defparam prom_inst_0.INIT_RAM_15 = 256'h99525E7559788B282BDABA5282452A7D2954A09BE2FA5EA9ABE17E8A2FA54B5D;
defparam prom_inst_0.INIT_RAM_16 = 256'hD2EEFABBCBCAA6BDD6DA75576D45C7E6EA5156D45A90749DE752D6E6179FBB5F;
defparam prom_inst_0.INIT_RAM_17 = 256'h9A18152796881BA3386CE4E4ECDD2D650141F66B532C88ABDB9472FC99A21C71;
defparam prom_inst_0.INIT_RAM_18 = 256'hB285153107CC85A5041B89E39D1717E1A529C8A518E5D26BC8912FF2B5B46D26;
defparam prom_inst_0.INIT_RAM_19 = 256'h14954174B495D78FC410835E5AF68505A76E3DFCB1C54A509E71C508374B2557;
defparam prom_inst_0.INIT_RAM_1A = 256'h5A4A16AEF5256276B4D564A6D4D6AC0EC48A5BC7AD259349C889978CE8D00336;
defparam prom_inst_0.INIT_RAM_1B = 256'hE889B8AE622C7FC2C56741DA5228D4C21721F2978BB956D5696D07B59285D498;
defparam prom_inst_0.INIT_RAM_1C = 256'h7D6FEAAAA01ECE9D974467B96A5644A3379B44C58067888CA484881C62D64D6A;
defparam prom_inst_0.INIT_RAM_1D = 256'h6E499C9A7EFE4D615E916E18AA14F2657AD624931E8C6D7C5B994B2AF7AA49DA;
defparam prom_inst_0.INIT_RAM_1E = 256'hF59DB1F88BAC76DE9C577E7072ACBD6FABF1FB5969FBF94D97BAD6D8A7B4A77D;
defparam prom_inst_0.INIT_RAM_1F = 256'hA7314BDA9169696D79795797A95AB01DFAEC75BBBCAAEFEDD246ED181D48D67A;
defparam prom_inst_0.INIT_RAM_20 = 256'h41CA1A7F4BD5B3825A6B8FC56CBAD8EE3B8A00852489D592CA7B3D6E375C7229;
defparam prom_inst_0.INIT_RAM_21 = 256'hB5418548965A4D6A86E6A86A09AAA28B2AEABA2C628626AC8B15B2D67B921B49;
defparam prom_inst_0.INIT_RAM_22 = 256'h163D8F5BD54961F74905E708E06195B91507057FE774B14A4D599C5F2593592D;
defparam prom_inst_0.INIT_RAM_23 = 256'h52931CB7DEFC9049A9FE1C6F4BE943C68B769955BBE955BA944957D63C82FB59;
defparam prom_inst_0.INIT_RAM_24 = 256'hD9FFEAE2EE6A85AD249185A45EE22AE897B1DD62E28898B1E226EC56FC8992E5;
defparam prom_inst_0.INIT_RAM_25 = 256'hEB6CA1DAD925524949A6A2B37D495F4954A1797EF6284B491A71556895E66145;
defparam prom_inst_0.INIT_RAM_26 = 256'hFE9EFFD796FDA12DAE767E7E57B57377E35D2D5BF5F34E41CCBA92476D2ABBB2;
defparam prom_inst_0.INIT_RAM_27 = 256'h296905BBDB4A55D14DCFDEACB54863D7B69597AD641DA52D57E455B5FA17EE6E;
defparam prom_inst_0.INIT_RAM_28 = 256'h61941C410E1E78BA73A14D255A5A5272C715B5454969ADA7BB2EEEC10534B374;
defparam prom_inst_0.INIT_RAM_29 = 256'hC3E8696129941F3A256869599259D05FF0A382A2B2F92B5BFF5D3561D06E4D7E;
defparam prom_inst_0.INIT_RAM_2A = 256'hD4A564B5E97A1DAD7D5FE5A1D2DA699875B756905E7955F2A57DE5A1DEF7B696;
defparam prom_inst_0.INIT_RAM_2B = 256'h8795172294985C9D254F135F5E4D12BDBB05555511E1D121790CEEF89456875B;
defparam prom_inst_0.INIT_RAM_2C = 256'hD4566BBCE85F5E5BE97D5621FBB595E79A17AD13B74859FE84EEFB4B736DB759;
defparam prom_inst_0.INIT_RAM_2D = 256'h7BBF3A173DB0A5A75A7929B9B93939B8C9752E561C1448BBD53524A89FF52DD6;
defparam prom_inst_0.INIT_RAM_2E = 256'h5F1CEE045C7B2938EE5E8C97929DB1C9F4BF7F24ED5D569D169CE7A64E7229E9;
defparam prom_inst_0.INIT_RAM_2F = 256'hDFC236FAFECCF05BE3389D91097951961E1CFE22DE321569DE9159E4A5245FE2;
defparam prom_inst_0.INIT_RAM_30 = 256'hD8326C62275E7DCFF9176FAFEFC080023D2B84DD03B9D3B402F7E55EF6223482;
defparam prom_inst_0.INIT_RAM_31 = 256'h979005EDA5521D56117975041749C49545D5443459D3B7624A46B400FCFFEF47;
defparam prom_inst_0.INIT_RAM_32 = 256'h56D465B21551BFF4AB2ACAB057BE756104185DB5787CFFEF5A75E527C96BE455;
defparam prom_inst_0.INIT_RAM_33 = 256'hD43F9A37BF0775FEA32DFCE7775F952C920F2755B3F695D5AE46C6F1F7EFF0B4;
defparam prom_inst_0.INIT_RAM_34 = 256'h119917545EC6FFDFFFFE6589FE245EEEE45DA44BA5DDA74B72991DFF2C8DD049;
defparam prom_inst_0.INIT_RAM_35 = 256'hAEE966E7E66DFE484057DD72B61229D70ED48213090ACE96D4FFD52F2B27235E;
defparam prom_inst_0.INIT_RAM_36 = 256'h3CAFFF75961ED5E49455D355451E05D85D76F0DE83FE8DB1671E9BAAFB1FFCDF;
defparam prom_inst_0.INIT_RAM_37 = 256'h29CBAC91556B3E2F85E61B4F4945DDDC5FBA7174978108B6E89D5545A4BD2617;
defparam prom_inst_0.INIT_RAM_38 = 256'h08030C6001E9E9F4157F3A2A8E360BB63992822B09C971E1C93BF9FAFB39B559;
defparam prom_inst_0.INIT_RAM_39 = 256'h5379257A8A9789E06D461054D580C4969C6956952ADE542FEC62875651617841;
defparam prom_inst_0.INIT_RAM_3A = 256'hCBA0594948575F7569415515697A141B549850103FEA08A2BB0200E416598795;
defparam prom_inst_0.INIT_RAM_3B = 256'h9E569855587DD61E691465247FFFBC9E44DEE834ACBE7B797F44218B8081A5FF;
defparam prom_inst_0.INIT_RAM_3C = 256'h5A5DB5C55546667A031D7D1878559877A53C362B9C05F7E981E6981DDF6ADDC6;
defparam prom_inst_0.INIT_RAM_3D = 256'hDC8235029549056FC914A5245CEE5250D2D2454AF9DC9D40E88C9C646436CA3E;
defparam prom_inst_0.INIT_RAM_3E = 256'h5241CE97D7B722B9282F8AF35573D4FBD0772E8AEFF32E8AECB55FFDC8210AD7;
defparam prom_inst_0.INIT_RAM_3F = 256'h08E548457F18830F3F5CC9E82F8AD7D7B8F752DBD072D57FF1F22BF00BF06165;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hBE30BAB63128C490C29B29B280A1D80A0D2C3098A8B8A838308C000800000010;
defparam prom_inst_1.INIT_RAM_01 = 256'hC3FCB400CC2C73FC8832C0362D8832C03E0C320030C800C01C00C8BFBFEC8DBE;
defparam prom_inst_1.INIT_RAM_02 = 256'h2B18B754AC6AB8EFBC30273C302B2CBCF4F98E30EEFFA39DBF1ACA708F4F3AE8;
defparam prom_inst_1.INIT_RAM_03 = 256'h3C32239CA3D8F0C883020C898B27F12E99B98B832F2D2D2CE62E3C3852B19555;
defparam prom_inst_1.INIT_RAM_04 = 256'h1E0E95A0681B06BE4281318082007000104104390C42FFF01E4FB3F01F2E2AF6;
defparam prom_inst_1.INIT_RAM_05 = 256'h70144F8F01F0C0002BC1DF0200F0C40C0BB7043480C3C1F0F080CC11A83A1783;
defparam prom_inst_1.INIT_RAM_06 = 256'h40D3402010CB304D2182FC10C7CB2FFC3CD0C03FDB4C41E49BD784F33FFFAE55;
defparam prom_inst_1.INIT_RAM_07 = 256'hBA61FD408DDD670C118E75DC208EEB8841801634802C300DC00B573C2DF3C146;
defparam prom_inst_1.INIT_RAM_08 = 256'h82608866232C7414200282D4416042B11762B17516F322F0A9C88CF028CC8035;
defparam prom_inst_1.INIT_RAM_09 = 256'hD4D11B4DD5D139538459CD7519BB59511831FB33F6378584262C348F70B5CC2C;
defparam prom_inst_1.INIT_RAM_0A = 256'h147F6603760575013C0712DF1E0511436FE59307BD406D6C5587DFD734D31504;
defparam prom_inst_1.INIT_RAM_0B = 256'hFE3EDC9A16D6615778664803144DDEC9594D31E0C25F70030E44101ED3F373EE;
defparam prom_inst_1.INIT_RAM_0C = 256'h34732BD710CF58D437DC5D31C51338E35A29EECBDE11DFDDEF537EE5AECC8DDD;
defparam prom_inst_1.INIT_RAM_0D = 256'h9130CE108402EC380C10BCC0000B000443C88D2D6F6EA827A127AA408D393F18;
defparam prom_inst_1.INIT_RAM_0E = 256'h976238E3E8FD73B12BB2C30C31C330A73E25EFF4DE84A58A8E305F5283239A88;
defparam prom_inst_1.INIT_RAM_0F = 256'h17601A6012108C086905F91A9D633358019DFD4BE34AF33C5D4EC4CE1DCE8FC3;
defparam prom_inst_1.INIT_RAM_10 = 256'h2282081A3C038C8E10473890EF4E23D30A4F4EB00A83C0493888EC4180000184;
defparam prom_inst_1.INIT_RAM_11 = 256'h82B7604B760B88FD68506EF98FBBFECD3A26E36E3C073332338FE394C2047C00;
defparam prom_inst_1.INIT_RAM_12 = 256'h39923E69E3B980434680002030BA89DB14CB2EA9C00AA2808ADB8F28E0BB9986;
defparam prom_inst_1.INIT_RAM_13 = 256'h30A87BA639005C0EC55B0EEBBBE6399F2F9ECE2784E33B91AEFEB13102CEE392;
defparam prom_inst_1.INIT_RAM_14 = 256'h13EDAEB4884C8D9C3FB1318FDDECC08FB989290A63518465888338C382E39234;
defparam prom_inst_1.INIT_RAM_15 = 256'h05E004DD3F21D010AA0B8F710A4012FC1960429A244A3DA3A1243DA2A1E30EB9;
defparam prom_inst_1.INIT_RAM_16 = 256'h8C93224C618AF32B110E454BEB4F8E03BE0052B4F670C390657BA2823190E669;
defparam prom_inst_1.INIT_RAM_17 = 256'h80DB74E3430433D98E343E32B6E8CBC2277FA63ABF388CBC94E421D61FE19823;
defparam prom_inst_1.INIT_RAM_18 = 256'h1A8E85230272E0AD00098C6DAF3E3BB8F822C4A6007E8C0A78DC641C60EC4C43;
defparam prom_inst_1.INIT_RAM_19 = 256'h339EFF47C3945CF08278A40C089C8E2065E6F38623BB79CD8E63BB9B028712AA;
defparam prom_inst_1.INIT_RAM_1A = 256'hCAC23393046720F300F4E59C3C3E32A7684E0C8104EC1C3071FE4F473EA259C2;
defparam prom_inst_1.INIT_RAM_1B = 256'hBDBDEAFA7BA8E9368FABC3A9F6BCFE0FFEABAA7DBDDF82762B174E5CF88CCE08;
defparam prom_inst_1.INIT_RAM_1C = 256'hDB70F0DF398A42E08F6C2238EE3F007892B419DBE6D29C9421918579F44E4F3E;
defparam prom_inst_1.INIT_RAM_1D = 256'hCD39F376672E2776DA75F010CF4E05F4104E2D043C4D4FC8CD18CDFC32BE64A9;
defparam prom_inst_1.INIT_RAM_1E = 256'h938D238E3F28E27278F84D26ED9F94EF8D63E939D99CB8278FFC4ECBF40F9F80;
defparam prom_inst_1.INIT_RAM_1F = 256'hEAC232FAF02B6F271B4BD4D9C4CC040C3C38E224C79D334772D4F6019E15F164;
defparam prom_inst_1.INIT_RAM_20 = 256'h4309A6317A33B1ED1331888C469A4C43184706E020075CD1A9D89CE53F78E0FC;
defparam prom_inst_1.INIT_RAM_21 = 256'h0E03AD083DA9CB315A73AD633BE6F1BDE3E8FAB8C1CCFE679E33300644CA384C;
defparam prom_inst_1.INIT_RAM_22 = 256'h08B22C2048336382330DDABEB6FBDA4E61201CC27E41A0F9CB18E8DD18BD3849;
defparam prom_inst_1.INIT_RAM_23 = 256'h4E7A38C07EFB30C3983D0FA3383B4EE1A212F7D44C36D33A9103436030A5DB38;
defparam prom_inst_1.INIT_RAM_24 = 256'h01000218018E8C68A8808CE848C29C82B2A3CCCC8503F0A3CEFCE8CCF6BF4CD4;
defparam prom_inst_1.INIT_RAM_25 = 256'h00B0A38AACA51330029C6FDE48375439811412200048C6220817492845062301;
defparam prom_inst_1.INIT_RAM_26 = 256'hD0800AAAC640231887DEA848C2AD40000224E01017C0360470CE62D104E304CB;
defparam prom_inst_1.INIT_RAM_27 = 256'h67A70CE690E9D744DF234A90430C2F30A29B6C24E808A82A280DC8AD22341313;
defparam prom_inst_1.INIT_RAM_28 = 256'h546D79C300B520D9DC7070E60C0000188E3C9D010908C0E74D6213031D7DC00D;
defparam prom_inst_1.INIT_RAM_29 = 256'h5033F8EBEF6D71CF3008EB30C408C6E8233626A69F3D0680014C7E1FD6D31F43;
defparam prom_inst_1.INIT_RAM_2A = 256'h28704419AF5A38A8613434A38A867188E0A01290003941DEB22007A32DF0A293;
defparam prom_inst_1.INIT_RAM_2B = 256'h7C7C5DEF519C307065722005C2DA21E9E69C254021230A230B64130C54128E1A;
defparam prom_inst_1.INIT_RAM_2C = 256'h4D73A4C367D12731D7448023AE60A0095230BA125E183700AFD30C1442134E09;
defparam prom_inst_1.INIT_RAM_2D = 256'h74C3B9F898F07D7029DFE76AFDD957E7091351F1FDBD8644107D325ADCD35002;
defparam prom_inst_1.INIT_RAM_2E = 256'hEA3B46FCF8DCE710C7E488F1FE74A38D6C46C43CC4E10A7A0272ED87EED07D06;
defparam prom_inst_1.INIT_RAM_2F = 256'h672AFB1B3B4EC9CD64B2F6046F19D2C23A3BD022469AB02F62FF207F9DCCF12C;
defparam prom_inst_1.INIT_RAM_30 = 256'hE60322E91BB6FB4F7C8BB1B33504CC4E0E1C6344AB144B97A4F96984DC39B5AC;
defparam prom_inst_1.INIT_RAM_31 = 256'h458800484AF3AF00802B1B000DE44E09D06D44404C4D9BCA440980081EF9EFAF;
defparam prom_inst_1.INIT_RAM_32 = 256'h80404B332F5137E08E3380E5BFDABC230108EC88B3DEF9EF86286609ED893116;
defparam prom_inst_1.INIT_RAM_33 = 256'hFB37C69194111B5619AB52C13BE99E2460AD3138994A04468084465AD96D98BF;
defparam prom_inst_1.INIT_RAM_34 = 256'h7AC4ABDA2E6BFD643DD712B10651213131284812BE90641A93C42F51104C4026;
defparam prom_inst_1.INIT_RAM_35 = 256'h2B89FA0CAA0A8A8E202176699F06BC4A32A2B18DEF2EB79EB677601A3A3A38AE;
defparam prom_inst_1.INIT_RAM_36 = 256'h0C5459808E3A00AC4AD5696CADAAB0932760A49ABF3819A31E381EEF8A3FD6FA;
defparam prom_inst_1.INIT_RAM_37 = 256'hF504DB1C13CDE8BAB01239F5FF72781BCB1AF803F7ADE84D806F48549E785D06;
defparam prom_inst_1.INIT_RAM_38 = 256'h0810841002906B11480409F25DFDF245E897F23EF9B300A32FE2BE1E3674AD59;
defparam prom_inst_1.INIT_RAM_39 = 256'h0ADB81A8463A2C69E82239C235AF31010F2B4235F2BD9625A70DABC2FF238A00;
defparam prom_inst_1.INIT_RAM_3A = 256'h45588BC8E88BFC1B6F2755B01BCE327AD608C0003FFA3868DF1729200DF4AD74;
defparam prom_inst_1.INIT_RAM_3B = 256'h85C238E708F82236F4908A92C1999086F77C9D10587FAADBB5F088C472A7BED4;
defparam prom_inst_1.INIT_RAM_3C = 256'hAD37F1427803631ABCEF83F8E8C338CB9711995D9C02ED3CA46F8A56F5F06F4F;
defparam prom_inst_1.INIT_RAM_3D = 256'h0023BFE388730E00333F9DCCF2311CE2313CCF809FC3E600EBF9CEEDE1F39CA6;
defparam prom_inst_1.INIT_RAM_3E = 256'h1CC371E076AB3AD5AE1C8E0B6ABB36CB3029152BDFFB152BD542047002390EFE;
defparam prom_inst_1.INIT_RAM_3F = 256'h0E238E05C030C020CF372ECE3D8E2076A4DF61DB70250811C1133226422A3912;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h8C327E343210C848F300100107E1307E13123CF0788078823CC40004000C0013;
defparam prom_inst_2.INIT_RAM_01 = 256'hCC3C88E20620030C4CB1333A214CB133322082B3320ACCC45C44FB0C30C0EC8C;
defparam prom_inst_2.INIT_RAM_02 = 256'h33DE6084CF6AA8CB0C408C8C408D70C08083EC3300C3D83D4F31C4320D8C13FE;
defparam prom_inst_2.INIT_RAM_03 = 256'h2080811C4360820208182062CCD4BB30AD5ACC2332323130490030C0133DC001;
defparam prom_inst_2.INIT_RAM_04 = 256'h238C630731CC73BEF39CFCF27204CC92CF3CF33420602A24AAA80324BA0021D8;
defparam prom_inst_2.INIT_RAM_05 = 256'hAFCAAAA24BA2AAAA90B9AA204206A4BA000AE9A2EBB81BA22432A38B1EB10013;
defparam prom_inst_2.INIT_RAM_06 = 256'hEAB9015BED00EFABEA803BBBAA8002AAAAB6AAAA80BABAAAE2AE2A8AAAAAC200;
defparam prom_inst_2.INIT_RAM_07 = 256'h7A0320023F8C0FB233204602EF700CCC1B7E8358FE412024C200BAE802AEAAEE;
defparam prom_inst_2.INIT_RAM_08 = 256'hEBFE8AEAFE02EEE6042F402BAEF210CDD8090981A9E7E5E7213276C4513184FC;
defparam prom_inst_2.INIT_RAM_09 = 256'h0114405104004054041410011D1D9D9DD711D5195599159BD51CEEFA800EBBA2;
defparam prom_inst_2.INIT_RAM_0A = 256'h4540061406050110004014101054451440041410001100010104101445045445;
defparam prom_inst_2.INIT_RAM_0B = 256'h0370302220240640809090101950101000110105050005545011541007F401AA;
defparam prom_inst_2.INIT_RAM_0C = 256'h483010041510438104100044145574DB6DF1331112CC66673445722723123013;
defparam prom_inst_2.INIT_RAM_0D = 256'hA880EF08AB0020AA3BCBBF000000000441C0405F539515511D9DD0C00C1E1E10;
defparam prom_inst_2.INIT_RAM_0E = 256'h98188208D23D08CFCC5049141141CBE105B8D7E5EC0328480C420830200480BE;
defparam prom_inst_2.INIT_RAM_0F = 256'h8482C84DCA88110728D303C533C8FE1074212323C8240CBE60A33F8D0EC813DC;
defparam prom_inst_2.INIT_RAM_10 = 256'hBC8CB2C8CBEDBEB2CAEEC831CEAE84ABA2EC3213B88BAA23BAA200DB75BBA7B2;
defparam prom_inst_2.INIT_RAM_11 = 256'h333B0FE8D8DF36FC080549F17F21FC8FDC4C0B08BF50DEF08B23CF8B2FF2ABAE;
defparam prom_inst_2.INIT_RAM_12 = 256'h88108C08C80033F3FF155D80462313C217730CCD164E2C3203616FA2043C2F5A;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFC133C5B10663670E421CC331C0301C03300CC3FF88323FC4F00FE0D8000810;
defparam prom_inst_2.INIT_RAM_14 = 256'h990000C13E223030082FEFC3E6060F7C0C00DCFC1BCD4FFC022BB1C700C81082;
defparam prom_inst_2.INIT_RAM_15 = 256'h1330BE3200FEC0FBE3210D8FBEB9F9BDF98BEFA00BD48E101F514D0C8BC8AD0A;
defparam prom_inst_2.INIT_RAM_16 = 256'hB2998CEE0303FF80C0BEBD261C902043BD4049C908452CABE880B4C84FAA6641;
defparam prom_inst_2.INIT_RAM_17 = 256'hB203BF23EF8CFFF48C747236744B28168C8880CA3FF22DFE8203A0006C111248;
defparam prom_inst_2.INIT_RAM_18 = 256'h81116E480610466205055F72D8408374F2F803E8FC60B2CA127F210C2B33FB2F;
defparam prom_inst_2.INIT_RAM_19 = 256'h4CA3083CECA8200C208208B6B28D102328D5D7A00880612336888020CA45DE66;
defparam prom_inst_2.INIT_RAM_1A = 256'h32144C99AB68851FAD4F7711000CB8CF0C032E284FF33ECA104F334105A8D368;
defparam prom_inst_2.INIT_RAM_1B = 256'hF22E32CCB002200D20C614A1043D430B200C20430CD8250890904241C513A151;
defparam prom_inst_2.INIT_RAM_1C = 256'h18C48D1141F73F1322CFFDE20C83D8C03DC8989807CDC303FDBDAD850CF79404;
defparam prom_inst_2.INIT_RAM_1D = 256'hFBCA32CC2F8904B62C4608FCEF50460A00FF03EFABAA9C8221022CC52DC0A7A1;
defparam prom_inst_2.INIT_RAM_1E = 256'hBFD008A32CC22909C20862A628D01FF02C4813DD30BE244423C4FF32F642100B;
defparam prom_inst_2.INIT_RAM_1F = 256'hEC4ACA31C4989C9094A61EDC033E401304322FA66107B8CCC02BAAAFCC980B40;
defparam prom_inst_2.INIT_RAM_20 = 256'h149DD39053FDD4D9FB73DC23E05E4D53574757F32C942011A104B37F500208BF;
defparam prom_inst_2.INIT_RAM_21 = 256'h409452C98D21144750B52D8B62DCB52C4160DC321ADD31D1248DE63E22158018;
defparam prom_inst_2.INIT_RAM_22 = 256'h6BCEB2712CC4DCA2C453B22CB4B2DAA0117661CA62ADA5211477F2000263DF6A;
defparam prom_inst_2.INIT_RAM_23 = 256'hC84089810B2C4518541C837370B15F91CF9DC63122B61DE62594D1F571F95DDD;
defparam prom_inst_2.INIT_RAM_24 = 256'hA62A9C9DC9DC132B27351325BF909D363FC8037DC964C64819315237204C37B1;
defparam prom_inst_2.INIT_RAM_25 = 256'h42F604B29F2E51DACA110BDEAB0016DA2D8ADCABB5810ECAB28482C8029C4445;
defparam prom_inst_2.INIT_RAM_26 = 256'h067BBA8A7E46043B220D60DCFA52EEC110377BFA882EC8C1115C5C0C4F76266F;
defparam prom_inst_2.INIT_RAM_27 = 256'hC4845266A42110C5144237413D851C7FAC98610F7C2B23282900F552544E999B;
defparam prom_inst_2.INIT_RAM_28 = 256'h106185145103FCE10452FB28B2B6B680224241DADADB2B2AAC4F999461514EE0;
defparam prom_inst_2.INIT_RAM_29 = 256'hDC0432015C6188453BA110DCF6EB953A88B6373733B2622EEBBA7054A5089CAB;
defparam prom_inst_2.INIT_RAM_2A = 256'h800BE6F2DC704B28414EB604B2B241C12EAEACA0BED843C45CEBE5448C2FACBC;
defparam prom_inst_2.INIT_RAM_2B = 256'h626150552DAD494B6862AEE13E0942AA223E41BC6A84A684F80F99ACC41812FA;
defparam prom_inst_2.INIT_RAM_2C = 256'h7143166885050FDD98143A04A22E8BE0404F855242D945110A88AE90A69452FA;
defparam prom_inst_2.INIT_RAM_2D = 256'hAAE941404DC43C42E1188452F42018E415584185494002A2A8700757E29840FE;
defparam prom_inst_2.INIT_RAM_2E = 256'h0C888F01021884FFB6052B818845088753C514E3B7004848E1C1614B1714BCB1;
defparam prom_inst_2.INIT_RAM_2F = 256'hF2A54797971984084E6506F6D8E535D1C98B915CF73D449C61C6856211110511;
defparam prom_inst_2.INIT_RAM_30 = 256'h81C051D10075D71AEF603939310C0045C22E13F6C4736631D70D78379CB1E914;
defparam prom_inst_2.INIT_RAM_31 = 256'h29E503ABBD82184B5318D8040716616404607D34CF62B60E0EC58004075D71CA;
defparam prom_inst_2.INIT_RAM_32 = 256'hE1FF3771F32CD4A3FEFFB3EF6380611C0486014243875D713BA7A99E4A73BDA9;
defparam prom_inst_2.INIT_RAM_33 = 256'h8316F73DC43D980503DC113BA60B51CC17E42DB53C462F698FF3731E1D75D7DF;
defparam prom_inst_2.INIT_RAM_34 = 256'h0FB6362798F2473E9F73D8409D0D48899D8B6ADA70AB6ADA32F6D87138336041;
defparam prom_inst_2.INIT_RAM_35 = 256'h0B43B18D51DA959CF08DC7F753777F603B495045D85DFA51C8D40A1E3E3E3E25;
defparam prom_inst_2.INIT_RAM_36 = 256'h87400D844184126375180D4F53094D73DCD34DE40167174840870D8B54825109;
defparam prom_inst_2.INIT_RAM_37 = 256'h2CBEB7077BCCD936F301C53514FDC73434B60D414E5E53EB6ED8B69A412A60A9;
defparam prom_inst_2.INIT_RAM_38 = 256'h00208908024AD8B5C2EEEC4448EB4EE35342DCFE70702E9C9046879797227184;
defparam prom_inst_2.INIT_RAM_39 = 256'h35145B4401044F762D31861181511DADA798D1017DCFC54C0DB536118698A580;
defparam prom_inst_2.INIT_RAM_3A = 256'hC083263A4F2610989C98B134C62D8987259600003FFA7AB0B8F606001416518D;
defparam prom_inst_2.INIT_RAM_3B = 256'hA6110610470501851AB5998E63BB43A714DC9FC8C8C27714004B30C0BCD87002;
defparam prom_inst_2.INIT_RAM_3C = 256'h069C7A690501D3DD74D8414726218600498B4685CC00171A5751A5FD8517D861;
defparam prom_inst_2.INIT_RAM_3D = 256'hBB2FD423F60450BB844211110438910F6F61103FD860C400EACEDCDCDFE3C8F4;
defparam prom_inst_2.INIT_RAM_3E = 256'h8114124908E374C4CDD52D76EA9D417540A0C033200CC03321CD8EEBB2FC8F53;
defparam prom_inst_2.INIT_RAM_3F = 256'h00080F2C8CFCC0008F9124FDF42D4908EF42ED5500A7363BB8B0F441F4423C4D;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0F003C3F33BCCEC0C0DCBDCBEFC1FEFC1F00303EF07EF070300700030003002F;
defparam prom_inst_3.INIT_RAM_01 = 256'hC7C03CC0C80C70C00B30C00C1C0B30C0001C310000C4002EE2EC00C30C3C0C0C;
defparam prom_inst_3.INIT_RAM_02 = 256'h033718CC0CC030F3CCB0300CB0359474343F0F31FC30C3E7303DCB73DDC72CF0;
defparam prom_inst_3.INIT_RAM_03 = 256'h0C3032DCB77C30C4C3230C4E43C3010C240243030D0D0D0C3F1F1C7E30335003;
defparam prom_inst_3.INIT_RAM_04 = 256'h1F2EFFEC0B02C0FCC0C0000000007030000000000C0000451555004515430DDF;
defparam prom_inst_3.INIT_RAM_05 = 256'h00105504515400001055154554540514500555045001515445FFC301BCFB80B0;
defparam prom_inst_3.INIT_RAM_06 = 256'h5451555155005545555005514550015454540015505551545455455000550055;
defparam prom_inst_3.INIT_RAM_07 = 256'hC31E1C33D91439003E2CB3C82041C7CB0108410FC8312C0C32C0555501555155;
defparam prom_inst_3.INIT_RAM_08 = 256'h50001055554100545540401545542C700F10BCF1365920F001C004F0F0C00F65;
defparam prom_inst_3.INIT_RAM_09 = 256'h7555DD7575D5D755D5D5D75CC884C44C440C444CCC848C0880CC545550055554;
defparam prom_inst_3.INIT_RAM_0A = 256'h575D5C5DDC5D755D5755D5D5D5755D7555D575D5755757575D5D5DD7575D55D5;
defparam prom_inst_3.INIT_RAM_0B = 256'h1333033385C55C571717175D7175D5757575D75D75D75D75D75D75D75EA75FAA;
defparam prom_inst_3.INIT_RAM_0C = 256'hC70D555555555415555555554514914D24510021030032220323002030032333;
defparam prom_inst_3.INIT_RAM_0D = 256'h711EC400554014141550BC030C32C00000CCE761EE682B672A242D00C135353C;
defparam prom_inst_3.INIT_RAM_0E = 256'h0F3032C340C110330700000000000041C3C43B1B30008C30C43FC33CF003C3E5;
defparam prom_inst_3.INIT_RAM_0F = 256'hC3CF203F214F0C008CFE0FCF0F8B12F2FD2F1F2C0B2CB03C3CC0CCB0B24B0FC0;
defparam prom_inst_3.INIT_RAM_10 = 256'h30320820B84104002046030F314543510C85400D1C32802E15C1C38100110DC8;
defparam prom_inst_3.INIT_RAM_11 = 256'h3EDD0F8D5CF73DD4C0CCC333CD0E0C36107873433400123C300C313C81085841;
defparam prom_inst_3.INIT_RAM_12 = 256'h302C34B0032C1CC08CC00007000E1E52DC40DC3300F7FD3F0E70DD02C3B50E0F;
defparam prom_inst_3.INIT_RAM_13 = 256'h1143074B32FF3C03C3F3CC731DCB72CC73C1CCF34C8302E30774732000B1C32C;
defparam prom_inst_3.INIT_RAM_14 = 256'h111F3CB2E4472F0FC7E3033372F3FC40781C113073FC38CC72F2DE790C032C30;
defparam prom_inst_3.INIT_RAM_15 = 256'hF3C0040FC7110730C2F3CCB30CFF31FC33FCC332CB80372C2E03172C7243C0BF;
defparam prom_inst_3.INIT_RAM_16 = 256'hC0D10F841E2CD10F38C4CFF3C3C32C70B560FC3C3830F03C4C30FCFC313044C0;
defparam prom_inst_3.INIT_RAM_17 = 256'h080C9C0FC13F33300F3F30303FFC803D43C7CF03C032CF34F4433041CC7BF10B;
defparam prom_inst_3.INIT_RAM_18 = 256'h470C8FCB001C371F0282EC81CF0CBC7DDF3040CF331FC0231C2482C7330CC881;
defparam prom_inst_3.INIT_RAM_19 = 256'h3030C7CE303F0C0F1071C7C4C0C30C008C3659F1CB07C0F2C4CB071C7F013C01;
defparam prom_inst_3.INIT_RAM_1A = 256'hC02C30110C8CB0C13C3C4E0C31C333B954003310B840E4031C2F3F31C31430CC;
defparam prom_inst_3.INIT_RAM_1B = 256'h31CF1EC7BC72C2CF2C33C320CFB432F31CB44832ED47FC7FC7C72F1F0B0C42F0;
defparam prom_inst_3.INIT_RAM_1C = 256'hC7CB0732C7844C1F0EF0C120C0300007E10FCF8F1E2100C4C20200B2C384C3CB;
defparam prom_inst_3.INIT_RAM_1D = 256'h4B233C03C90FCBC3F032CF300D1CB3C8C7840155154550F2F2C0C10B810BEF00;
defparam prom_inst_3.INIT_RAM_1E = 256'hE130CB32CC72CC7CF2C7F132C001D841CD4B1E130F243FCB0C0B840CDF0C0C3C;
defparam prom_inst_3.INIT_RAM_1F = 256'h4C75033C3BC7C3C7CBF0FC7C73C40C00CBB2F13441C210B83015551553CF22CF;
defparam prom_inst_3.INIT_RAM_20 = 256'hC33940183D811CFB111E432C41DA0C731EC10DDC820B0C3000C7E8430CF2C734;
defparam prom_inst_3.INIT_RAM_21 = 256'h0FC30F2034C0C30EC3B3ECB33ECF32EC702DC372C0CF0CF1C0B120C4C45435C0;
defparam prom_inst_3.INIT_RAM_22 = 256'h8E5B961CC7C7C3FFC70FBCEF333ECD4423333C3F1FF230C0C30CD2F40F0E108F;
defparam prom_inst_3.INIT_RAM_23 = 256'hC03CB03CF14470C340EFB83C2C2032B379DC30FF4410F121F303FC921F944410;
defparam prom_inst_3.INIT_RAM_24 = 256'hF1C00B2472470C8C80C80C85C48F3473C10B6040330C30CB430C32C461C344BC;
defparam prom_inst_3.INIT_RAM_25 = 256'h0C90C3C8C08F3013200CF353FFC7F713F20C23F11CB0C02148C3F3200FCBC303;
defparam prom_inst_3.INIT_RAM_26 = 256'h52F110C34441C30080C335C33F3FC44C70104110034447C01C07835C7843C449;
defparam prom_inst_3.INIT_RAM_27 = 256'h83030F44F0C0FC01C73E440E1101659130030CF8400C8C8CC0B5333F0C3F11C1;
defparam prom_inst_3.INIT_RAM_28 = 256'hC80CB2C30C361220C70F900FC8C8C8C72C0F1F2323208C8D447911C33F1CB475;
defparam prom_inst_3.INIT_RAM_29 = 256'h8F0730CC030CB070DC40C710081042DCCB32E2E2E13340F441C43FC372D1CFC1;
defparam prom_inst_3.INIT_RAM_2A = 256'h001C41E3432C3C8F1CB811C3C8C82C00F1313030041303870FF040C30C41303C;
defparam prom_inst_3.INIT_RAM_2B = 256'h0F0F2C70B2343CBC8F0C5470C451404344E7FFFFD7C3FD43117B1106F2070F13;
defparam prom_inst_3.INIT_RAM_2C = 256'h1CB0C44071F3391183CCC4C304413C411C31117F1F2030C0305107CFF0030F13;
defparam prom_inst_3.INIT_RAM_2D = 256'hD4410C7DDA5C2323C0C7033CF31C0372E3C33C3C34B501443F3F012E77833F44;
defparam prom_inst_3.INIT_RAM_2E = 256'hF4B0791C32C70320C1F1E8FC7031CB031CB1CF3CC1F7F03F7CF02C3300C337D4;
defparam prom_inst_3.INIT_RAM_2F = 256'h9651D919196832C0700C73C887D1FCFC3C3C0F8388E43F032C31331C0F1C33C1;
defparam prom_inst_3.INIT_RAM_30 = 256'h4C7054730D965966448D919191F2333036B4478870D880E5436510C88FF35543;
defparam prom_inst_3.INIT_RAM_31 = 256'h0CC5008C84B0CFF10807CB0280C82C81CF2FDE320481E3E264E18802D1451472;
defparam prom_inst_3.INIT_RAM_32 = 256'h7F3CC1C32DF315B484210C402F073FC30200F55F0D11451488F08C35030E123C;
defparam prom_inst_3.INIT_RAM_33 = 256'hFCE0C8E207C20B473E431C3EC3F11C36CF61A213E471F08C7A4C0C44451440C0;
defparam prom_inst_3.INIT_RAM_34 = 256'hBD88D3F30F9E10140101231C04023111123C85230FFC8F23DB48CF3C80148020;
defparam prom_inst_3.INIT_RAM_35 = 256'h330F3CF030FCC303903CF1D82DC8B48CC93C701C47A0B61C3F957FE4E4E4E4E0;
defparam prom_inst_3.INIT_RAM_36 = 256'h34E204BF0C30FF1CF3FF65F33FFC3F0CC3C71E70C1A0C1CB1CB0DC331CB45430;
defparam prom_inst_3.INIT_RAM_37 = 256'hC00003C13C010F33CB0032C2C7CC32F1F3E1DC907E0F1C002C0FC8CC0E2F3CCC;
defparam prom_inst_3.INIT_RAM_38 = 256'h0010C02A033F87324F44431CC0001C041F1CC3340C3CC7C3070C191919030FF1;
defparam prom_inst_3.INIT_RAM_39 = 256'hF3CB233CECF3EC83E08033FCBF0CB23231C7FCFF2C377C3878B3D3FC3103F000;
defparam prom_inst_3.INIT_RAM_3A = 256'h40ECC0CC3CC3C7CBC3CFFFCFC0C43CF0FCC0E02817DA52D8515843DC01C00CBF;
defparam prom_inst_3.INIT_RAM_3B = 256'h02FCF0C7F0CC9032C05C6E592D111CC3C04BB432121750CB1A30C8C0C30F0C68;
defparam prom_inst_3.INIT_RAM_3C = 256'h3003132075807B2032CF1CF0F0FCF0E4E9E06863840930C00F2C00F8F2C30F2C;
defparam prom_inst_3.INIT_RAM_3D = 256'h1103430348C70FD1C70C0F1C33D1F1F37371C3CC473C3F80695B6752614F644D;
defparam prom_inst_3.INIT_RAM_3E = 256'h31C31C3CFD7C3CCC0F31CC318000701C703D3303300533033472346110340D0D;
defparam prom_inst_3.INIT_RAM_3F = 256'h01C3C2EDCB30030CBF31C30F33CC3CFD7C3D833CF031C8D1B0130330C3303402;

endmodule //Gowin_pROM
