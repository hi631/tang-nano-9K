//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.03
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Fri Nov 25 17:28:28 2022

module Gowin_pROM_boot (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire [15:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h1E89C806C8041F0E5152550E16539090A3C404A390C3B9D2505612348EE0D28C;
defparam prom_inst_0.INIT_RAM_01 = 256'h19E8E800C80E03F0EBE8E8C803F478E8A103048104A1BCD08ED88CFC02A38B36;
defparam prom_inst_0.INIT_RAM_02 = 256'h495358435841E246E804048AB903070E368BE8CF02C41F025D5F595B06260416;
defparam prom_inst_0.INIT_RAM_03 = 256'h03DD8B26E83A04328A46E81846043C048EC8C0B410B953435053535353445042;
defparam prom_inst_0.INIT_RAM_04 = 256'hF300C90000BE03FA74020A74800F5A01C17F67E8F0E2C300C3D257E80AF94303;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFBD000204B9BF000000F300000000BECA2010BEBBA415B9BFC02AEBBFC9C900;
defparam prom_inst_0.INIT_RAM_06 = 256'h287501658AC802B80176048ABE0203954BBE068EE8C5036E38064BE80E8C468A;
defparam prom_inst_0.INIT_RAM_07 = 256'h805133E873FC7573EB01057568EBE86D2FE874FCEBFE567834B8E8C000BC756E;
defparam prom_inst_0.INIT_RAM_08 = 256'h087514EBE8194FE8E8213AE8133C1375801D3C35BFE8693C00F47566EB010575;
defparam prom_inst_0.INIT_RAM_09 = 256'hBAE704E88AC8EF02C28BB702B7C3E800D10373FC02168BFFC3000475C3D27400;
defparam prom_inst_0.INIT_RAM_0A = 256'h05758017CBE8E8E00B7580FFC3A500B9BFE0C3078926B80826C0C08E8B00C3EF;
defparam prom_inst_0.INIT_RAM_0B = 256'h05B9C2E9B80036016E016DC3E8FF0AE814E8E809C3E25BBA097645E802FAEB09;
defparam prom_inst_0.INIT_RAM_0C = 256'hC30700BA0DFC8AC8C3EF8B015208E4E86FFCAAF3ABF300FC8B01CA8BE8FAC3A5;
defparam prom_inst_0.INIT_RAM_0D = 256'h8B26E846892600FE00FCEB5E0DFC742E248ABE00560101948A26E8F274748AC8;
defparam prom_inst_0.INIT_RAM_0E = 256'hA3E874E08A2626C80204F9808B3FB0C88900C83400D4301630BBBFEB88260159;
defparam prom_inst_0.INIT_RAM_0F = 256'h8B50E850E03826C80204F9800E8B3E8B0146B0CF36065801C48AE8015800F78B;
defparam prom_inst_0.INIT_RAM_10 = 256'h04B5C30000EEB0000F2400B103C2E8C1C300C810D2E2060200D88A0000E0001C;
defparam prom_inst_0.INIT_RAM_11 = 256'hE846F7EB75208A0000BAC358E80DC358E820C3E5FE00F1754200009C048AB1FF;
defparam prom_inst_0.INIT_RAM_12 = 256'h3C0000B4B0E0302C2437724072305859D00AC15A1689F000520CFE04F980FF3C;
defparam prom_inst_0.INIT_RAM_13 = 256'h30040272C358E80F0008E8C0C3005800C48AE075C4FE8800ECEB4E00F474800D;
defparam prom_inst_0.INIT_RAM_14 = 256'hE80684045AEEBA58C084EC035052EC03F9748024FDBAE2FFBAFD08758024FFBA;
defparam prom_inst_0.INIT_RAM_15 = 256'h000000000000000000000000000000000000000000000000003E36386D0DEB46;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'hE858E8F8C28BDA830010E0C1C1D074C03BE8E80100BEAAE8E9CCD08ED88EFCFA;
defparam prom_inst_0.INIT_RAM_31 = 256'hEB8340009EE8E8007474023E7565003EE8E2C38183011F755949E851DB331FE8;
defparam prom_inst_0.INIT_RAM_32 = 256'h33FF00EAA5F3100033E0A4F3B9FBB4BE01008EE4754B8800DC8AE8FCA7E8BEF9;
defparam prom_inst_0.INIT_RAM_33 = 256'hFF330068B042B04AB042B04AB042B003EE0810B0BA06E6403243B08FB08BB080;
defparam prom_inst_0.INIT_RAM_34 = 256'h40E402E8FA52DABAC307C084F7FE01B4BEFF8EB806C3EE2AEE0103C8ABF3B80C;
defparam prom_inst_0.INIT_RAM_35 = 256'h06B9E8C34725E7E8E2FFACC39090909001B4C3F8E4E8E40A81F5D002EC0040E4;
defparam prom_inst_0.INIT_RAM_36 = 256'h9BE8E8FBB50EFC80E8160A06FFD6054401B4BAF451B28A5074FF0574D3E8FFE7;
defparam prom_inst_0.INIT_RAM_37 = 256'hB8BEAAFC58FFFC8B04B1CCFEE8CE6575FF9EA0BEB4FB87E8B903C3FFEFC0FF98;
defparam prom_inst_0.INIT_RAM_38 = 256'h31E8E12B117580FF1975FF4FACBE5840FF528BE1B1FFCEBE74CC71E8BEFFFF77;
defparam prom_inst_0.INIT_RAM_39 = 256'h6F20697477204B387361647244536F20657370206E2049428BFFEFC08B41F64D;
defparam prom_inst_0.INIT_RAM_3A = 256'hFF0000770000FF0000490100950000402E2E30303030202C6230353120325352;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000F000EA000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[15:0],dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 16;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hC80EDC8B2689168C505356571E0654C3C8068BC8D08C9ABC8E5878BBB8D000B8;
defparam prom_inst_1.INIT_RAM_01 = 256'h8E01001D5BE81E8BE803046F02A1E804C806FDE8E8C8CBC08EC08EC8FAC81A47;
defparam prom_inst_1.INIT_RAM_02 = 256'h494458445842C3F503AA39E8000479E8C80203C65C5B8307C4835E5A58C88BC8;
defparam prom_inst_1.INIT_RAM_03 = 256'h59E8E807042CB046E8040438EB4675208AC004A1BE0046535049202053452020;
defparam prom_inst_1.INIT_RAM_04 = 256'hBBA415B9BFC02C74801BFA8001FAE28048E8BA010974805201E8E20303758043;
defparam prom_inst_1.INIT_RAM_05 = 256'h2ECFE3FFE800002010BEBBA415B9BFC014EBBFCACA00F300CA0000BEC92010BE;
defparam prom_inst_1.INIT_RAM_06 = 256'hFC80643C8A0510BFE846663CC81172E8E8C5C838039F44BEE8C88E01C838C300;
defparam prom_inst_1.INIT_RAM_07 = 256'h70FCEB01057580143C5F51E86D3C0256EBFF0575807740E8BB12009D15BAE814;
defparam prom_inst_1.INIT_RAM_08 = 256'hFE80673C006EEB000039EB000575C68B70FC7562EB0005753EEBE8053C4716E8;
defparam prom_inst_1.INIT_RAM_09 = 256'h02F28A5BC0C438A1F0BA5300EB80001E08E8027580C88BCA47E904E8743CFF02;
defparam prom_inst_1.INIT_RAM_0A = 256'h4FE801FAEBFFFFB55BBA62FCF1E8F310E00000BE0A44F000448923B806F000B8;
defparam prom_inst_1.INIT_RAM_0B = 256'hF300FF33BE07680138016F01FF9A80E8E80009F8E4E8FFE005EBE80908758012;
defparam prom_inst_1.INIT_RAM_0C = 256'h11BF52F00375802411BE5AC241E8EB09057480C302EB047480C25DE801628BFC;
defparam prom_inst_1.INIT_RAM_0D = 256'hE80400A246141074805EE81C03758027FC80C810BEE805E8E80400D28B453C05;
defparam prom_inst_1.INIT_RAM_0E = 256'h500050173825058836067500044F8B003616CDE81689E8C889C8C35E4614CEEB;
defparam prom_inst_1.INIT_RAM_0F = 256'hE8F700661774258A36067500C834C83000B0E82EE2C8024715E8008E1DE859E8;
defparam prom_inst_1.INIT_RAM_10 = 256'hDDE8F28B21E8E83AC5E8C68BE8C28C04C68B9BE8BEC3C8364758E8C451E8E858;
defparam prom_inst_1.INIT_RAM_11 = 256'h0023048A46033C04B100515000BCB05000C4B05075CD0DE8C9FE0DE8E8462610;
defparam prom_inst_1.INIT_RAM_12 = 256'h750856E8C3FF8AC3C30F2C053C0C3CC3DAEB04E2C838C28EE281EBC174041C74;
defparam prom_inst_1.INIT_RAM_13 = 256'h24EB07040A3C00022458E804505001E805E850C30D3C460453E8CCFE5BE800FC;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFE474C08AC303FCF9758024FEBAC35AFCBAC084EC0352C3E05B8DE8003CEC03;
defparam prom_inst_1.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000000000000000D006E6FC3F4;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_30 = 256'hF89BF81EA2E85000C12BB90A06EA8B4E85F8F8BFB1E8E800F57400BCC08EC88C;
defparam prom_inst_1.INIT_RAM_31 = 256'h7540078ABB000060EB317800810A4E0081C3020000D2C083585A01445250C3F8;
defparam prom_inst_1.INIT_RAM_32 = 256'hE7C0FF009090E3FFB9F600BF00098BCCF000EAD433F746249DE800A28A000100;
defparam prom_inst_1.INIT_RAM_33 = 256'h00B907B8EE00EE0DEE00EE0CEE20EE0AD4BAB0EE03C0C340E6C0E634E70FE70B;
defparam prom_inst_1.INIT_RAM_34 = 256'hE802FA72C0ECB90380B4F775ACABE8ACCE5033C000B8EEEEB04201B8BA07012E;
defparam prom_inst_1.INIT_RAM_35 = 256'hE800FFDEF8E288FFC3FAEFE8ED90909090EEFFB0754038405BE973DCE8C008E8;
defparam prom_inst_1.INIT_RAM_36 = 256'hE8FFFFB48B0275FEFFD275E4C483E8FFC6EF03DA8B5250C2C3F5FC8046FFF633;
defparam prom_inst_1.INIT_RAM_37 = 256'hE8CE4B7580587BE8E12B5B75FF91A6BECCFEE8CEEF01E2FF000ADABA91E83341;
defparam prom_inst_1.INIT_RAM_38 = 256'h8BFFFC8B12B1FEFC51E8E40AE8CE2374A858E8FC2B0464E8BEEDFEFFCEB255E8;
defparam prom_inst_1.INIT_RAM_39 = 256'h206E676E69612C4220746C206143206E746E6572746F534FC3C10DE833E7CD86;
defparam prom_inst_1.INIT_RAM_3A = 256'h007A0000FF004069000087AA00480000002E2029313A30667370303231283332;
defparam prom_inst_1.INIT_RAM_3B = 256'h000000000000000000000000000000000000000000000000000000000000FF00;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h00000000000000CC000000000000000000000000000000000000000000000000;

endmodule //Gowin_pROM_boot
